import lynxTypes::*;

module crc32_calc(
    // Networking interface - Incoming and outgoing traffic 
    AXI4S.m m_axis_rx, 
    AXI4S.m m_axis_tx, 

    // Incoming clock and reset
    input logic nclk, 
    input logic nresetn
);

// Regs for the first pipeline stage 
logic stage_1_valid; 
logic [511:0] stage_1_data;
logic [511:0] stage_1_masked_data; 
logic [63:0] stage_1_keep;
logic stage_1_last; 
logic [7:0] ai_word_count; 

// Regs for the second pipeline stage
logic stage_2_valid;
logic [511:0] stage_2_data_bypass; 
logic [31:0] stage_2_crc_value; 
logic [63:0] stage_2_keep; 
logic stage_2_last; 

// Calculation Factors for bitwise CRC 
logic [511:0] d; 
logic [31:0] c;

// Regs for the third pipeline stage 
logic stage_3_valid; 
logic [511:0] stage_3_data;
logic [63:0] stage_3_keep; 
logic stage_3_last; 
logic stall_pipeline; 
logic [31:0] stage_3_crc_value; 

// Regs for the fourth pipeline stage 
logic stage_4_valid; 
logic [511:0] stage_4_data; 
logic [63:0] stage_4_keep; 
logic stage_4_last; 
logic switch_output; 

// Bitmask for CRC-calculation 
logic [511:0] bitmask; 

// Parameter for the header length
param logic []


/////////////////////////////////////////////////////////////////////////////////////////////
//
// Assignment of d for CRC-calculation to stage_1_bitmasked data
//
/////////////////////////////////////////////////////////////////////////////////////////////
assign d = stage_1_bitmasked; 
assign c = stage_2_crc_value;   

always_ff @(posedge nclk) begin
    if(nresetn == 1'b0) begin 
        // Flush the pipeline: Reset the stage registers to 0
        stage_1_valid <= 1'b0;
        stage_1_data <= 512'b0;
        stage_1_keep <= 64'b0;
        stage_1_last <= 1'b0;
        stage_1_masked_data <= 512'b0;

        stage_2_valid <= 1'b0; 
        stage_2_data_bypass <= 512'b0;
        stage_2_keep <= 64'b0; 
        stage_2_last <= 1'b0; 
        stage_2_crc_value <= 32'b0; 

        stage_3_valid <= 1'b0; 
        stage_3_data <= 512'b0;
        stage_3_keep <= 64'b0;
        stage_3_last <= 1'b0;
        stall_pipeline <= 1'b0;
        stage_3_crc_value <= 32'b0;  

        stage_4_valid <= 1'b0; 
        stage_4_data <= 512'b0; 
        stage_4_keep <= 63'b0; 
        stage_4_last <= 1'b0;
        switch_output <= 1'b0; 

        // Set the required bits of the bitmask for the masking operation in this stage 
        bitmask[3:0] <= 4'b1; // Traffic Class
        bitmask[11:8] <= 4'b1; // Traffic Class
        bitmask[31:12] <= 20'b1; // Flow Label
        bitmask[63:56] <= 8'b1; // Hop Limit
        bitmask[383:56] <= 16'b1; // UDP checksum
        bitmask[423:416] <= 8'b1; // BTH Resv8a

        // Reset the CRC-seed to all 1
        stage_2_crc_value <= 32'b1;

        // Reset the ai word count 
        ai_word_count <= 0; 
    end 

    /////////////////////////////////////////////////////////////////////
    //
    // STAGE 1: LOADING AND BITMASKING
    //
    /////////////////////////////////////////////////////////////////////
    
    // Forward direct signals: valid, last, keep, data 
    stage_1_valid <= m_axis_rx.valid;
    stage_1_last <= m_axis_rx.last;
    stage_1_keep <= m_axis_rx.keep;
    stage_1_data <= m_axis_rx.data;

    // If input is valid, load and mask data - else it's just 0s 
    if(m_axis_rx.valid) begin 
        // Only mask the first word (only one with Header Fields)
        if(ai_word_count == 0) begin 
            stage_1_masked_data[423:0] <= m_axis_rx.data[423:0] | bitmask[423:0];
            stage_1_masked_data[511:424] <= m_axis_rx.data[511:424];

            // Reset the crc-seed value to all 1 for beginning of processing in the next step 
            stage_2_crc_value <= 32'b1; 
        end else begin
            stage_1_masked_data <= m_axis_rx.data;
        end 

        // Increment the ai_word_count if .last is not set 
        if(!m_axis_rx.last) begin
            ai_word_count <= ai_word_count + 1;
        end else begin 
            ai_word_count <= 0;
        end
    end


    ///////////////////////////////////////////////////////////////////////
    //
    // STAGE 2: CRC calculation
    //
    ///////////////////////////////////////////////////////////////////////

    // Forward direct signals: valid, last, keep, data
    stage_2_valid <= stage_1_valid; 
    stage_2_last <= stage_1_last; 
    stage_2_keep <= stage_1_keep;
    stage_2_data_bypass <= stage_1_data; 

    // Bitwise calculation of the CRC-value based on the bitmasked data and the CRC-seed. 
    stage_2_crc_value[0] = d[511] ^ d[510] ^ d[508] ^ d[507] ^ d[506] ^ d[502] ^ d[501] ^ d[500] ^ d[495] ^ d[494] ^ d[493] ^ d[492] ^ d[491] ^ d[490] ^ d[489] ^ d[488] ^ d[486] ^ d[483] ^ d[482] ^ d[481] ^ d[480] ^ d[479] ^ d[477] ^ d[476] ^ d[472] ^ d[470] ^ d[468] ^ d[465] ^ d[464] ^ d[462] ^ d[461] ^ d[458] ^ d[452] ^ d[450] ^ d[449] ^ d[448] ^ d[444] ^ d[437] ^ d[436] ^ d[434] ^ d[433] ^ d[424] ^ d[422] ^ d[419] ^ d[418] ^ d[416] ^ d[414] ^ d[412] ^ d[409] ^ d[408] ^ d[407] ^ d[405] ^ d[404] ^ d[400] ^ d[399] ^ d[398] ^ d[396] ^ d[393] ^ d[392] ^ d[391] ^ d[390] ^ d[388] ^ d[387] ^ d[386] ^ d[381] ^ d[378] ^ d[376] ^ d[374] ^ d[372] ^ d[369] ^ d[368] ^ d[366] ^ d[363] ^ d[362] ^ d[359] ^ d[358] ^ d[357] ^ d[353] ^ d[349] ^ d[348] ^ d[347] ^ d[345] ^ d[344] ^ d[342] ^ d[341] ^ d[339] ^ d[338] ^ d[337] ^ d[335] ^ d[334] ^ d[333] ^ d[328] ^ d[327] ^ d[322] ^ d[321] ^ d[320] ^ d[319] ^ d[318] ^ d[317] ^ d[315] ^ d[312] ^ d[310] ^ d[309] ^ d[305] ^ d[303] ^ d[302] ^ d[300] ^ d[299] ^ d[298] ^ d[297] ^ d[296] ^ d[295] ^ d[294] ^ d[292] ^ d[290] ^ d[288] ^ d[287] ^ d[286] ^ d[283] ^ d[279] ^ d[277] ^ d[276] ^ d[274] ^ d[273] ^ d[269] ^ d[268] ^ d[265] ^ d[264] ^ d[261] ^ d[259] ^ d[257] ^ d[255] ^ d[252] ^ d[248] ^ d[243] ^ d[237] ^ d[234] ^ d[230] ^ d[228] ^ d[227] ^ d[226] ^ d[224] ^ d[216] ^ d[214] ^ d[212] ^ d[210] ^ d[209] ^ d[208] ^ d[207] ^ d[203] ^ d[202] ^ d[201] ^ d[199] ^ d[198] ^ d[197] ^ d[194] ^ d[193] ^ d[192] ^ d[191] ^ d[190] ^ d[188] ^ d[186] ^ d[183] ^ d[182] ^ d[172] ^ d[171] ^ d[170] ^ d[169] ^ d[167] ^ d[166] ^ d[162] ^ d[161] ^ d[158] ^ d[156] ^ d[155] ^ d[151] ^ d[149] ^ d[144] ^ d[143] ^ d[137] ^ d[136] ^ d[135] ^ d[134] ^ d[132] ^ d[128] ^ d[127] ^ d[126] ^ d[125] ^ d[123] ^ d[119] ^ d[118] ^ d[117] ^ d[116] ^ d[114] ^ d[113] ^ d[111] ^ d[110] ^ d[106] ^ d[104] ^ d[103] ^ d[101] ^ d[99] ^ d[98] ^ d[97] ^ d[96] ^ d[95] ^ d[94] ^ d[87] ^ d[85] ^ d[84] ^ d[83] ^ d[82] ^ d[81] ^ d[79] ^ d[73] ^ d[72] ^ d[68] ^ d[67] ^ d[66] ^ d[65] ^ d[63] ^ d[61] ^ d[60] ^ d[58] ^ d[55] ^ d[54] ^ d[53] ^ d[50] ^ d[48] ^ d[47] ^ d[45] ^ d[44] ^ d[37] ^ d[34] ^ d[32] ^ d[31] ^ d[30] ^ d[29] ^ d[28] ^ d[26] ^ d[25] ^ d[24] ^ d[16] ^ d[12] ^ d[10] ^ d[9] ^ d[6] ^ d[0] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[6] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[15] ^ c[20] ^ c[21] ^ c[22] ^ c[26] ^ c[27] ^ c[28] ^ c[30] ^ c[31];
    stage_2_crc_value[1] = d[510] ^ d[509] ^ d[506] ^ d[503] ^ d[500] ^ d[496] ^ d[488] ^ d[487] ^ d[486] ^ d[484] ^ d[479] ^ d[478] ^ d[476] ^ d[473] ^ d[472] ^ d[471] ^ d[470] ^ d[469] ^ d[468] ^ d[466] ^ d[464] ^ d[463] ^ d[461] ^ d[459] ^ d[458] ^ d[453] ^ d[452] ^ d[451] ^ d[448] ^ d[445] ^ d[444] ^ d[438] ^ d[436] ^ d[435] ^ d[433] ^ d[425] ^ d[424] ^ d[423] ^ d[422] ^ d[420] ^ d[418] ^ d[417] ^ d[416] ^ d[415] ^ d[414] ^ d[413] ^ d[412] ^ d[410] ^ d[407] ^ d[406] ^ d[404] ^ d[401] ^ d[398] ^ d[397] ^ d[396] ^ d[394] ^ d[390] ^ d[389] ^ d[386] ^ d[382] ^ d[381] ^ d[379] ^ d[378] ^ d[377] ^ d[376] ^ d[375] ^ d[374] ^ d[373] ^ d[372] ^ d[370] ^ d[368] ^ d[367] ^ d[366] ^ d[364] ^ d[362] ^ d[360] ^ d[357] ^ d[354] ^ d[353] ^ d[350] ^ d[347] ^ d[346] ^ d[344] ^ d[343] ^ d[341] ^ d[340] ^ d[337] ^ d[336] ^ d[333] ^ d[329] ^ d[327] ^ d[323] ^ d[317] ^ d[316] ^ d[315] ^ d[313] ^ d[312] ^ d[311] ^ d[309] ^ d[306] ^ d[305] ^ d[304] ^ d[302] ^ d[301] ^ d[294] ^ d[293] ^ d[292] ^ d[291] ^ d[290] ^ d[289] ^ d[286] ^ d[284] ^ d[283] ^ d[280] ^ d[279] ^ d[278] ^ d[276] ^ d[275] ^ d[273] ^ d[270] ^ d[268] ^ d[266] ^ d[264] ^ d[262] ^ d[261] ^ d[260] ^ d[259] ^ d[258] ^ d[257] ^ d[256] ^ d[255] ^ d[253] ^ d[252] ^ d[249] ^ d[248] ^ d[244] ^ d[243] ^ d[238] ^ d[237] ^ d[235] ^ d[234] ^ d[231] ^ d[230] ^ d[229] ^ d[226] ^ d[225] ^ d[224] ^ d[217] ^ d[216] ^ d[215] ^ d[214] ^ d[213] ^ d[212] ^ d[211] ^ d[207] ^ d[204] ^ d[201] ^ d[200] ^ d[197] ^ d[195] ^ d[190] ^ d[189] ^ d[188] ^ d[187] ^ d[186] ^ d[184] ^ d[182] ^ d[173] ^ d[169] ^ d[168] ^ d[166] ^ d[163] ^ d[161] ^ d[159] ^ d[158] ^ d[157] ^ d[155] ^ d[152] ^ d[151] ^ d[150] ^ d[149] ^ d[145] ^ d[143] ^ d[138] ^ d[134] ^ d[133] ^ d[132] ^ d[129] ^ d[125] ^ d[124] ^ d[123] ^ d[120] ^ d[116] ^ d[115] ^ d[113] ^ d[112] ^ d[110] ^ d[107] ^ d[106] ^ d[105] ^ d[103] ^ d[102] ^ d[101] ^ d[100] ^ d[94] ^ d[88] ^ d[87] ^ d[86] ^ d[81] ^ d[80] ^ d[79] ^ d[74] ^ d[72] ^ d[69] ^ d[65] ^ d[64] ^ d[63] ^ d[62] ^ d[60] ^ d[59] ^ d[58] ^ d[56] ^ d[53] ^ d[51] ^ d[50] ^ d[49] ^ d[47] ^ d[46] ^ d[44] ^ d[38] ^ d[37] ^ d[35] ^ d[34] ^ d[33] ^ d[28] ^ d[27] ^ d[24] ^ d[17] ^ d[16] ^ d[13] ^ d[12] ^ d[11] ^ d[9] ^ d[7] ^ d[6] ^ d[1] ^ d[0] ^ c[4] ^ c[6] ^ c[7] ^ c[8] ^ c[16] ^ c[20] ^ c[23] ^ c[26] ^ c[29] ^ c[30];
    stage_2_crc_value[2] = d[508] ^ d[506] ^ d[504] ^ d[502] ^ d[500] ^ d[497] ^ d[495] ^ d[494] ^ d[493] ^ d[492] ^ d[491] ^ d[490] ^ d[487] ^ d[486] ^ d[485] ^ d[483] ^ d[482] ^ d[481] ^ d[476] ^ d[474] ^ d[473] ^ d[471] ^ d[469] ^ d[468] ^ d[467] ^ d[461] ^ d[460] ^ d[459] ^ d[458] ^ d[454] ^ d[453] ^ d[450] ^ d[448] ^ d[446] ^ d[445] ^ d[444] ^ d[439] ^ d[433] ^ d[426] ^ d[425] ^ d[423] ^ d[422] ^ d[421] ^ d[417] ^ d[415] ^ d[413] ^ d[412] ^ d[411] ^ d[409] ^ d[404] ^ d[402] ^ d[400] ^ d[397] ^ d[396] ^ d[395] ^ d[393] ^ d[392] ^ d[388] ^ d[386] ^ d[383] ^ d[382] ^ d[381] ^ d[380] ^ d[379] ^ d[377] ^ d[375] ^ d[373] ^ d[372] ^ d[371] ^ d[367] ^ d[366] ^ d[365] ^ d[362] ^ d[361] ^ d[359] ^ d[357] ^ d[355] ^ d[354] ^ d[353] ^ d[351] ^ d[349] ^ d[339] ^ d[335] ^ d[333] ^ d[330] ^ d[327] ^ d[324] ^ d[322] ^ d[321] ^ d[320] ^ d[319] ^ d[316] ^ d[315] ^ d[314] ^ d[313] ^ d[309] ^ d[307] ^ d[306] ^ d[300] ^ d[299] ^ d[298] ^ d[297] ^ d[296] ^ d[293] ^ d[291] ^ d[288] ^ d[286] ^ d[285] ^ d[284] ^ d[283] ^ d[281] ^ d[280] ^ d[273] ^ d[271] ^ d[268] ^ d[267] ^ d[264] ^ d[263] ^ d[262] ^ d[260] ^ d[258] ^ d[256] ^ d[255] ^ d[254] ^ d[253] ^ d[252] ^ d[250] ^ d[249] ^ d[248] ^ d[245] ^ d[244] ^ d[243] ^ d[239] ^ d[238] ^ d[237] ^ d[236] ^ d[235] ^ d[234] ^ d[232] ^ d[231] ^ d[228] ^ d[225] ^ d[224] ^ d[218] ^ d[217] ^ d[215] ^ d[213] ^ d[210] ^ d[209] ^ d[207] ^ d[205] ^ d[203] ^ d[199] ^ d[197] ^ d[196] ^ d[194] ^ d[193] ^ d[192] ^ d[189] ^ d[187] ^ d[186] ^ d[185] ^ d[182] ^ d[174] ^ d[172] ^ d[171] ^ d[166] ^ d[164] ^ d[161] ^ d[160] ^ d[159] ^ d[155] ^ d[153] ^ d[152] ^ d[150] ^ d[149] ^ d[146] ^ d[143] ^ d[139] ^ d[137] ^ d[136] ^ d[133] ^ d[132] ^ d[130] ^ d[128] ^ d[127] ^ d[124] ^ d[123] ^ d[121] ^ d[119] ^ d[118] ^ d[110] ^ d[108] ^ d[107] ^ d[102] ^ d[99] ^ d[98] ^ d[97] ^ d[96] ^ d[94] ^ d[89] ^ d[88] ^ d[85] ^ d[84] ^ d[83] ^ d[80] ^ d[79] ^ d[75] ^ d[72] ^ d[70] ^ d[68] ^ d[67] ^ d[64] ^ d[59] ^ d[58] ^ d[57] ^ d[55] ^ d[53] ^ d[52] ^ d[51] ^ d[44] ^ d[39] ^ d[38] ^ d[37] ^ d[36] ^ d[35] ^ d[32] ^ d[31] ^ d[30] ^ d[26] ^ d[24] ^ d[18] ^ d[17] ^ d[16] ^ d[14] ^ d[13] ^ d[9] ^ d[8] ^ d[7] ^ d[6] ^ d[2] ^ d[1] ^ d[0] ^ c[1] ^ c[2] ^ c[3] ^ c[5] ^ c[6] ^ c[7] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[15] ^ c[17] ^ c[20] ^ c[22] ^ c[24] ^ c[26] ^ c[28];
    stage_2_crc_value[3] = d[509] ^ d[507] ^ d[505] ^ d[503] ^ d[501] ^ d[498] ^ d[496] ^ d[495] ^ d[494] ^ d[493] ^ d[492] ^ d[491] ^ d[488] ^ d[487] ^ d[486] ^ d[484] ^ d[483] ^ d[482] ^ d[477] ^ d[475] ^ d[474] ^ d[472] ^ d[470] ^ d[469] ^ d[468] ^ d[462] ^ d[461] ^ d[460] ^ d[459] ^ d[455] ^ d[454] ^ d[451] ^ d[449] ^ d[447] ^ d[446] ^ d[445] ^ d[440] ^ d[434] ^ d[427] ^ d[426] ^ d[424] ^ d[423] ^ d[422] ^ d[418] ^ d[416] ^ d[414] ^ d[413] ^ d[412] ^ d[410] ^ d[405] ^ d[403] ^ d[401] ^ d[398] ^ d[397] ^ d[396] ^ d[394] ^ d[393] ^ d[389] ^ d[387] ^ d[384] ^ d[383] ^ d[382] ^ d[381] ^ d[380] ^ d[378] ^ d[376] ^ d[374] ^ d[373] ^ d[372] ^ d[368] ^ d[367] ^ d[366] ^ d[363] ^ d[362] ^ d[360] ^ d[358] ^ d[356] ^ d[355] ^ d[354] ^ d[352] ^ d[350] ^ d[340] ^ d[336] ^ d[334] ^ d[331] ^ d[328] ^ d[325] ^ d[323] ^ d[322] ^ d[321] ^ d[320] ^ d[317] ^ d[316] ^ d[315] ^ d[314] ^ d[310] ^ d[308] ^ d[307] ^ d[301] ^ d[300] ^ d[299] ^ d[298] ^ d[297] ^ d[294] ^ d[292] ^ d[289] ^ d[287] ^ d[286] ^ d[285] ^ d[284] ^ d[282] ^ d[281] ^ d[274] ^ d[272] ^ d[269] ^ d[268] ^ d[265] ^ d[264] ^ d[263] ^ d[261] ^ d[259] ^ d[257] ^ d[256] ^ d[255] ^ d[254] ^ d[253] ^ d[251] ^ d[250] ^ d[249] ^ d[246] ^ d[245] ^ d[244] ^ d[240] ^ d[239] ^ d[238] ^ d[237] ^ d[236] ^ d[235] ^ d[233] ^ d[232] ^ d[229] ^ d[226] ^ d[225] ^ d[219] ^ d[218] ^ d[216] ^ d[214] ^ d[211] ^ d[210] ^ d[208] ^ d[206] ^ d[204] ^ d[200] ^ d[198] ^ d[197] ^ d[195] ^ d[194] ^ d[193] ^ d[190] ^ d[188] ^ d[187] ^ d[186] ^ d[183] ^ d[175] ^ d[173] ^ d[172] ^ d[167] ^ d[165] ^ d[162] ^ d[161] ^ d[160] ^ d[156] ^ d[154] ^ d[153] ^ d[151] ^ d[150] ^ d[147] ^ d[144] ^ d[140] ^ d[138] ^ d[137] ^ d[134] ^ d[133] ^ d[131] ^ d[129] ^ d[128] ^ d[125] ^ d[124] ^ d[122] ^ d[120] ^ d[119] ^ d[111] ^ d[109] ^ d[108] ^ d[103] ^ d[100] ^ d[99] ^ d[98] ^ d[97] ^ d[95] ^ d[90] ^ d[89] ^ d[86] ^ d[85] ^ d[84] ^ d[81] ^ d[80] ^ d[76] ^ d[73] ^ d[71] ^ d[69] ^ d[68] ^ d[65] ^ d[60] ^ d[59] ^ d[58] ^ d[56] ^ d[54] ^ d[53] ^ d[52] ^ d[45] ^ d[40] ^ d[39] ^ d[38] ^ d[37] ^ d[36] ^ d[33] ^ d[32] ^ d[31] ^ d[27] ^ d[25] ^ d[19] ^ d[18] ^ d[17] ^ d[15] ^ d[14] ^ d[10] ^ d[9] ^ d[8] ^ d[7] ^ d[3] ^ d[2] ^ d[1] ^ c[2] ^ c[3] ^ c[4] ^ c[6] ^ c[7] ^ c[8] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[15] ^ c[16] ^ c[18] ^ c[21] ^ c[23] ^ c[25] ^ c[27] ^ c[29];
    stage_2_crc_value[4] = d[511] ^ d[507] ^ d[504] ^ d[501] ^ d[500] ^ d[499] ^ d[497] ^ d[496] ^ d[491] ^ d[490] ^ d[487] ^ d[486] ^ d[485] ^ d[484] ^ d[482] ^ d[481] ^ d[480] ^ d[479] ^ d[478] ^ d[477] ^ d[475] ^ d[473] ^ d[472] ^ d[471] ^ d[469] ^ d[468] ^ d[465] ^ d[464] ^ d[463] ^ d[460] ^ d[458] ^ d[456] ^ d[455] ^ d[449] ^ d[447] ^ d[446] ^ d[444] ^ d[441] ^ d[437] ^ d[436] ^ d[435] ^ d[434] ^ d[433] ^ d[428] ^ d[427] ^ d[425] ^ d[423] ^ d[422] ^ d[418] ^ d[417] ^ d[416] ^ d[415] ^ d[413] ^ d[412] ^ d[411] ^ d[409] ^ d[408] ^ d[407] ^ d[406] ^ d[405] ^ d[402] ^ d[400] ^ d[397] ^ d[396] ^ d[395] ^ d[394] ^ d[393] ^ d[392] ^ d[391] ^ d[387] ^ d[386] ^ d[385] ^ d[384] ^ d[383] ^ d[382] ^ d[379] ^ d[378] ^ d[377] ^ d[376] ^ d[375] ^ d[373] ^ d[372] ^ d[367] ^ d[366] ^ d[364] ^ d[362] ^ d[361] ^ d[358] ^ d[356] ^ d[355] ^ d[351] ^ d[349] ^ d[348] ^ d[347] ^ d[345] ^ d[344] ^ d[342] ^ d[339] ^ d[338] ^ d[334] ^ d[333] ^ d[332] ^ d[329] ^ d[328] ^ d[327] ^ d[326] ^ d[324] ^ d[323] ^ d[320] ^ d[319] ^ d[316] ^ d[312] ^ d[311] ^ d[310] ^ d[308] ^ d[305] ^ d[303] ^ d[301] ^ d[297] ^ d[296] ^ d[294] ^ d[293] ^ d[292] ^ d[285] ^ d[282] ^ d[279] ^ d[277] ^ d[276] ^ d[275] ^ d[274] ^ d[270] ^ d[268] ^ d[266] ^ d[262] ^ d[261] ^ d[260] ^ d[259] ^ d[258] ^ d[256] ^ d[254] ^ d[251] ^ d[250] ^ d[248] ^ d[247] ^ d[246] ^ d[245] ^ d[243] ^ d[241] ^ d[240] ^ d[239] ^ d[238] ^ d[236] ^ d[233] ^ d[228] ^ d[224] ^ d[220] ^ d[219] ^ d[217] ^ d[216] ^ d[215] ^ d[214] ^ d[211] ^ d[210] ^ d[208] ^ d[205] ^ d[203] ^ d[202] ^ d[197] ^ d[196] ^ d[195] ^ d[193] ^ d[192] ^ d[190] ^ d[189] ^ d[187] ^ d[186] ^ d[184] ^ d[183] ^ d[182] ^ d[176] ^ d[174] ^ d[173] ^ d[172] ^ d[171] ^ d[170] ^ d[169] ^ d[168] ^ d[167] ^ d[163] ^ d[158] ^ d[157] ^ d[156] ^ d[154] ^ d[152] ^ d[149] ^ d[148] ^ d[145] ^ d[144] ^ d[143] ^ d[141] ^ d[139] ^ d[138] ^ d[137] ^ d[136] ^ d[130] ^ d[129] ^ d[128] ^ d[127] ^ d[121] ^ d[120] ^ d[119] ^ d[118] ^ d[117] ^ d[116] ^ d[114] ^ d[113] ^ d[112] ^ d[111] ^ d[109] ^ d[106] ^ d[103] ^ d[100] ^ d[97] ^ d[95] ^ d[94] ^ d[91] ^ d[90] ^ d[86] ^ d[84] ^ d[83] ^ d[79] ^ d[77] ^ d[74] ^ d[73] ^ d[70] ^ d[69] ^ d[68] ^ d[67] ^ d[65] ^ d[63] ^ d[59] ^ d[58] ^ d[57] ^ d[50] ^ d[48] ^ d[47] ^ d[46] ^ d[45] ^ d[44] ^ d[41] ^ d[40] ^ d[39] ^ d[38] ^ d[33] ^ d[31] ^ d[30] ^ d[29] ^ d[25] ^ d[24] ^ d[20] ^ d[19] ^ d[18] ^ d[15] ^ d[12] ^ d[11] ^ d[8] ^ d[6] ^ d[4] ^ d[3] ^ d[2] ^ d[0] ^ c[0] ^ c[1] ^ c[2] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[10] ^ c[11] ^ c[16] ^ c[17] ^ c[19] ^ c[20] ^ c[21] ^ c[24] ^ c[27] ^ c[31];
    stage_2_crc_value[5] = d[511] ^ d[510] ^ d[507] ^ d[506] ^ d[505] ^ d[498] ^ d[497] ^ d[495] ^ d[494] ^ d[493] ^ d[490] ^ d[489] ^ d[487] ^ d[485] ^ d[478] ^ d[477] ^ d[474] ^ d[473] ^ d[469] ^ d[468] ^ d[466] ^ d[462] ^ d[459] ^ d[458] ^ d[457] ^ d[456] ^ d[452] ^ d[449] ^ d[447] ^ d[445] ^ d[444] ^ d[442] ^ d[438] ^ d[435] ^ d[433] ^ d[429] ^ d[428] ^ d[426] ^ d[423] ^ d[422] ^ d[417] ^ d[413] ^ d[410] ^ d[406] ^ d[405] ^ d[404] ^ d[403] ^ d[401] ^ d[400] ^ d[399] ^ d[397] ^ d[395] ^ d[394] ^ d[391] ^ d[390] ^ d[385] ^ d[384] ^ d[383] ^ d[381] ^ d[380] ^ d[379] ^ d[377] ^ d[373] ^ d[372] ^ d[369] ^ d[367] ^ d[366] ^ d[365] ^ d[358] ^ d[356] ^ d[353] ^ d[352] ^ d[350] ^ d[347] ^ d[346] ^ d[344] ^ d[343] ^ d[342] ^ d[341] ^ d[340] ^ d[338] ^ d[337] ^ d[330] ^ d[329] ^ d[325] ^ d[324] ^ d[322] ^ d[319] ^ d[318] ^ d[315] ^ d[313] ^ d[311] ^ d[310] ^ d[306] ^ d[305] ^ d[304] ^ d[303] ^ d[300] ^ d[299] ^ d[296] ^ d[293] ^ d[292] ^ d[290] ^ d[288] ^ d[287] ^ d[280] ^ d[279] ^ d[278] ^ d[275] ^ d[274] ^ d[273] ^ d[271] ^ d[268] ^ d[267] ^ d[265] ^ d[264] ^ d[263] ^ d[262] ^ d[260] ^ d[251] ^ d[249] ^ d[247] ^ d[246] ^ d[244] ^ d[243] ^ d[242] ^ d[241] ^ d[240] ^ d[239] ^ d[230] ^ d[229] ^ d[228] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[221] ^ d[220] ^ d[218] ^ d[217] ^ d[215] ^ d[214] ^ d[211] ^ d[210] ^ d[208] ^ d[207] ^ d[206] ^ d[204] ^ d[202] ^ d[201] ^ d[199] ^ d[196] ^ d[192] ^ d[187] ^ d[186] ^ d[185] ^ d[184] ^ d[182] ^ d[177] ^ d[175] ^ d[174] ^ d[173] ^ d[168] ^ d[167] ^ d[166] ^ d[164] ^ d[162] ^ d[161] ^ d[159] ^ d[157] ^ d[156] ^ d[153] ^ d[151] ^ d[150] ^ d[146] ^ d[145] ^ d[143] ^ d[142] ^ d[140] ^ d[139] ^ d[138] ^ d[136] ^ d[135] ^ d[134] ^ d[132] ^ d[131] ^ d[130] ^ d[129] ^ d[127] ^ d[126] ^ d[125] ^ d[123] ^ d[122] ^ d[121] ^ d[120] ^ d[116] ^ d[115] ^ d[112] ^ d[111] ^ d[107] ^ d[106] ^ d[103] ^ d[99] ^ d[97] ^ d[94] ^ d[92] ^ d[91] ^ d[83] ^ d[82] ^ d[81] ^ d[80] ^ d[79] ^ d[78] ^ d[75] ^ d[74] ^ d[73] ^ d[72] ^ d[71] ^ d[70] ^ d[69] ^ d[67] ^ d[65] ^ d[64] ^ d[63] ^ d[61] ^ d[59] ^ d[55] ^ d[54] ^ d[53] ^ d[51] ^ d[50] ^ d[49] ^ d[46] ^ d[44] ^ d[42] ^ d[41] ^ d[40] ^ d[39] ^ d[37] ^ d[29] ^ d[28] ^ d[24] ^ d[21] ^ d[20] ^ d[19] ^ d[13] ^ d[10] ^ d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[3] ^ d[1] ^ d[0] ^ c[5] ^ c[7] ^ c[9] ^ c[10] ^ c[13] ^ c[14] ^ c[15] ^ c[17] ^ c[18] ^ c[25] ^ c[26] ^ c[27] ^ c[30] ^ c[31];
    stage_2_crc_value[6] = d[511] ^ d[508] ^ d[507] ^ d[506] ^ d[499] ^ d[498] ^ d[496] ^ d[495] ^ d[494] ^ d[491] ^ d[490] ^ d[488] ^ d[486] ^ d[479] ^ d[478] ^ d[475] ^ d[474] ^ d[470] ^ d[469] ^ d[467] ^ d[463] ^ d[460] ^ d[459] ^ d[458] ^ d[457] ^ d[453] ^ d[450] ^ d[448] ^ d[446] ^ d[445] ^ d[443] ^ d[439] ^ d[436] ^ d[434] ^ d[430] ^ d[429] ^ d[427] ^ d[424] ^ d[423] ^ d[418] ^ d[414] ^ d[411] ^ d[407] ^ d[406] ^ d[405] ^ d[404] ^ d[402] ^ d[401] ^ d[400] ^ d[398] ^ d[396] ^ d[395] ^ d[392] ^ d[391] ^ d[386] ^ d[385] ^ d[384] ^ d[382] ^ d[381] ^ d[380] ^ d[378] ^ d[374] ^ d[373] ^ d[370] ^ d[368] ^ d[367] ^ d[366] ^ d[359] ^ d[357] ^ d[354] ^ d[353] ^ d[351] ^ d[348] ^ d[347] ^ d[345] ^ d[344] ^ d[343] ^ d[342] ^ d[341] ^ d[339] ^ d[338] ^ d[331] ^ d[330] ^ d[326] ^ d[325] ^ d[323] ^ d[320] ^ d[319] ^ d[316] ^ d[314] ^ d[312] ^ d[311] ^ d[307] ^ d[306] ^ d[305] ^ d[304] ^ d[301] ^ d[300] ^ d[297] ^ d[294] ^ d[293] ^ d[291] ^ d[289] ^ d[288] ^ d[281] ^ d[280] ^ d[279] ^ d[276] ^ d[275] ^ d[274] ^ d[272] ^ d[269] ^ d[268] ^ d[266] ^ d[265] ^ d[264] ^ d[263] ^ d[261] ^ d[252] ^ d[250] ^ d[248] ^ d[247] ^ d[245] ^ d[244] ^ d[243] ^ d[242] ^ d[241] ^ d[240] ^ d[231] ^ d[230] ^ d[229] ^ d[228] ^ d[227] ^ d[226] ^ d[225] ^ d[222] ^ d[221] ^ d[219] ^ d[218] ^ d[216] ^ d[215] ^ d[212] ^ d[211] ^ d[209] ^ d[208] ^ d[207] ^ d[205] ^ d[203] ^ d[202] ^ d[200] ^ d[197] ^ d[193] ^ d[188] ^ d[187] ^ d[186] ^ d[185] ^ d[183] ^ d[178] ^ d[176] ^ d[175] ^ d[174] ^ d[169] ^ d[168] ^ d[167] ^ d[165] ^ d[163] ^ d[162] ^ d[160] ^ d[158] ^ d[157] ^ d[154] ^ d[152] ^ d[151] ^ d[147] ^ d[146] ^ d[144] ^ d[143] ^ d[141] ^ d[140] ^ d[139] ^ d[137] ^ d[136] ^ d[135] ^ d[133] ^ d[132] ^ d[131] ^ d[130] ^ d[128] ^ d[127] ^ d[126] ^ d[124] ^ d[123] ^ d[122] ^ d[121] ^ d[117] ^ d[116] ^ d[113] ^ d[112] ^ d[108] ^ d[107] ^ d[104] ^ d[100] ^ d[98] ^ d[95] ^ d[93] ^ d[92] ^ d[84] ^ d[83] ^ d[82] ^ d[81] ^ d[80] ^ d[79] ^ d[76] ^ d[75] ^ d[74] ^ d[73] ^ d[72] ^ d[71] ^ d[70] ^ d[68] ^ d[66] ^ d[65] ^ d[64] ^ d[62] ^ d[60] ^ d[56] ^ d[55] ^ d[54] ^ d[52] ^ d[51] ^ d[50] ^ d[47] ^ d[45] ^ d[43] ^ d[42] ^ d[41] ^ d[40] ^ d[38] ^ d[30] ^ d[29] ^ d[25] ^ d[22] ^ d[21] ^ d[20] ^ d[14] ^ d[11] ^ d[8] ^ d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[2] ^ d[1] ^ c[6] ^ c[8] ^ c[10] ^ c[11] ^ c[14] ^ c[15] ^ c[16] ^ c[18] ^ c[19] ^ c[26] ^ c[27] ^ c[28] ^ c[31];
    stage_2_crc_value[7] = d[511] ^ d[510] ^ d[509] ^ d[506] ^ d[502] ^ d[501] ^ d[499] ^ d[497] ^ d[496] ^ d[494] ^ d[493] ^ d[490] ^ d[488] ^ d[487] ^ d[486] ^ d[483] ^ d[482] ^ d[481] ^ d[477] ^ d[475] ^ d[472] ^ d[471] ^ d[465] ^ d[462] ^ d[460] ^ d[459] ^ d[454] ^ d[452] ^ d[451] ^ d[450] ^ d[448] ^ d[447] ^ d[446] ^ d[440] ^ d[436] ^ d[435] ^ d[434] ^ d[433] ^ d[431] ^ d[430] ^ d[428] ^ d[425] ^ d[422] ^ d[418] ^ d[416] ^ d[415] ^ d[414] ^ d[409] ^ d[406] ^ d[404] ^ d[403] ^ d[402] ^ d[401] ^ d[400] ^ d[398] ^ d[397] ^ d[391] ^ d[390] ^ d[388] ^ d[385] ^ d[383] ^ d[382] ^ d[379] ^ d[378] ^ d[376] ^ d[375] ^ d[372] ^ d[371] ^ d[367] ^ d[366] ^ d[363] ^ d[362] ^ d[360] ^ d[359] ^ d[357] ^ d[355] ^ d[354] ^ d[353] ^ d[352] ^ d[347] ^ d[346] ^ d[343] ^ d[341] ^ d[340] ^ d[338] ^ d[337] ^ d[335] ^ d[334] ^ d[333] ^ d[332] ^ d[331] ^ d[328] ^ d[326] ^ d[324] ^ d[322] ^ d[319] ^ d[318] ^ d[313] ^ d[310] ^ d[309] ^ d[308] ^ d[307] ^ d[306] ^ d[303] ^ d[301] ^ d[300] ^ d[299] ^ d[297] ^ d[296] ^ d[289] ^ d[288] ^ d[287] ^ d[286] ^ d[283] ^ d[282] ^ d[281] ^ d[280] ^ d[279] ^ d[275] ^ d[274] ^ d[270] ^ d[268] ^ d[267] ^ d[266] ^ d[262] ^ d[261] ^ d[259] ^ d[257] ^ d[255] ^ d[253] ^ d[252] ^ d[251] ^ d[249] ^ d[246] ^ d[245] ^ d[244] ^ d[242] ^ d[241] ^ d[237] ^ d[234] ^ d[232] ^ d[231] ^ d[229] ^ d[224] ^ d[223] ^ d[222] ^ d[220] ^ d[219] ^ d[217] ^ d[214] ^ d[213] ^ d[207] ^ d[206] ^ d[204] ^ d[202] ^ d[199] ^ d[197] ^ d[193] ^ d[192] ^ d[191] ^ d[190] ^ d[189] ^ d[187] ^ d[184] ^ d[183] ^ d[182] ^ d[179] ^ d[177] ^ d[176] ^ d[175] ^ d[172] ^ d[171] ^ d[168] ^ d[167] ^ d[164] ^ d[163] ^ d[162] ^ d[159] ^ d[156] ^ d[153] ^ d[152] ^ d[151] ^ d[149] ^ d[148] ^ d[147] ^ d[145] ^ d[143] ^ d[142] ^ d[141] ^ d[140] ^ d[138] ^ d[135] ^ d[133] ^ d[131] ^ d[129] ^ d[126] ^ d[124] ^ d[122] ^ d[119] ^ d[116] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[106] ^ d[105] ^ d[104] ^ d[103] ^ d[98] ^ d[97] ^ d[95] ^ d[93] ^ d[87] ^ d[80] ^ d[79] ^ d[77] ^ d[76] ^ d[75] ^ d[74] ^ d[71] ^ d[69] ^ d[68] ^ d[60] ^ d[58] ^ d[57] ^ d[56] ^ d[54] ^ d[52] ^ d[51] ^ d[50] ^ d[47] ^ d[46] ^ d[45] ^ d[43] ^ d[42] ^ d[41] ^ d[39] ^ d[37] ^ d[34] ^ d[32] ^ d[29] ^ d[28] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[16] ^ d[15] ^ d[10] ^ d[8] ^ d[7] ^ d[5] ^ d[3] ^ d[2] ^ d[0] ^ c[1] ^ c[2] ^ c[3] ^ c[6] ^ c[7] ^ c[8] ^ c[10] ^ c[13] ^ c[14] ^ c[16] ^ c[17] ^ c[19] ^ c[21] ^ c[22] ^ c[26] ^ c[29] ^ c[30] ^ c[31];
    stage_2_crc_value[8] = d[508] ^ d[506] ^ d[503] ^ d[501] ^ d[498] ^ d[497] ^ d[493] ^ d[492] ^ d[490] ^ d[487] ^ d[486] ^ d[484] ^ d[481] ^ d[480] ^ d[479] ^ d[478] ^ d[477] ^ d[473] ^ d[470] ^ d[468] ^ d[466] ^ d[465] ^ d[464] ^ d[463] ^ d[462] ^ d[460] ^ d[458] ^ d[455] ^ d[453] ^ d[451] ^ d[450] ^ d[447] ^ d[444] ^ d[441] ^ d[435] ^ d[433] ^ d[432] ^ d[431] ^ d[429] ^ d[426] ^ d[424] ^ d[423] ^ d[422] ^ d[418] ^ d[417] ^ d[415] ^ d[414] ^ d[412] ^ d[410] ^ d[409] ^ d[408] ^ d[403] ^ d[402] ^ d[401] ^ d[400] ^ d[396] ^ d[393] ^ d[390] ^ d[389] ^ d[388] ^ d[387] ^ d[384] ^ d[383] ^ d[381] ^ d[380] ^ d[379] ^ d[378] ^ d[377] ^ d[374] ^ d[373] ^ d[369] ^ d[367] ^ d[366] ^ d[364] ^ d[362] ^ d[361] ^ d[360] ^ d[359] ^ d[357] ^ d[356] ^ d[355] ^ d[354] ^ d[349] ^ d[345] ^ d[337] ^ d[336] ^ d[332] ^ d[329] ^ d[328] ^ d[325] ^ d[323] ^ d[322] ^ d[321] ^ d[318] ^ d[317] ^ d[315] ^ d[314] ^ d[312] ^ d[311] ^ d[308] ^ d[307] ^ d[305] ^ d[304] ^ d[303] ^ d[301] ^ d[299] ^ d[296] ^ d[295] ^ d[294] ^ d[292] ^ d[289] ^ d[286] ^ d[284] ^ d[282] ^ d[281] ^ d[280] ^ d[279] ^ d[277] ^ d[275] ^ d[274] ^ d[273] ^ d[271] ^ d[267] ^ d[265] ^ d[264] ^ d[263] ^ d[262] ^ d[261] ^ d[260] ^ d[259] ^ d[258] ^ d[257] ^ d[256] ^ d[255] ^ d[254] ^ d[253] ^ d[250] ^ d[248] ^ d[247] ^ d[246] ^ d[245] ^ d[242] ^ d[238] ^ d[237] ^ d[235] ^ d[234] ^ d[233] ^ d[232] ^ d[228] ^ d[227] ^ d[226] ^ d[225] ^ d[223] ^ d[221] ^ d[220] ^ d[218] ^ d[216] ^ d[215] ^ d[212] ^ d[210] ^ d[209] ^ d[205] ^ d[202] ^ d[201] ^ d[200] ^ d[199] ^ d[197] ^ d[186] ^ d[185] ^ d[184] ^ d[182] ^ d[180] ^ d[178] ^ d[177] ^ d[176] ^ d[173] ^ d[171] ^ d[170] ^ d[168] ^ d[167] ^ d[166] ^ d[165] ^ d[164] ^ d[163] ^ d[162] ^ d[161] ^ d[160] ^ d[158] ^ d[157] ^ d[156] ^ d[155] ^ d[154] ^ d[153] ^ d[152] ^ d[151] ^ d[150] ^ d[148] ^ d[146] ^ d[142] ^ d[141] ^ d[139] ^ d[137] ^ d[135] ^ d[130] ^ d[128] ^ d[126] ^ d[120] ^ d[119] ^ d[118] ^ d[116] ^ d[114] ^ d[113] ^ d[112] ^ d[109] ^ d[107] ^ d[105] ^ d[103] ^ d[101] ^ d[97] ^ d[95] ^ d[88] ^ d[87] ^ d[85] ^ d[84] ^ d[83] ^ d[82] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[76] ^ d[75] ^ d[73] ^ d[70] ^ d[69] ^ d[68] ^ d[67] ^ d[66] ^ d[65] ^ d[63] ^ d[60] ^ d[59] ^ d[57] ^ d[54] ^ d[52] ^ d[51] ^ d[50] ^ d[46] ^ d[45] ^ d[43] ^ d[42] ^ d[40] ^ d[38] ^ d[37] ^ d[35] ^ d[34] ^ d[33] ^ d[32] ^ d[31] ^ d[28] ^ d[23] ^ d[22] ^ d[17] ^ d[12] ^ d[11] ^ d[10] ^ d[8] ^ d[4] ^ d[3] ^ d[1] ^ d[0] ^ c[0] ^ c[1] ^ c[4] ^ c[6] ^ c[7] ^ c[10] ^ c[12] ^ c[13] ^ c[17] ^ c[18] ^ c[21] ^ c[23] ^ c[26] ^ c[28];
    stage_2_crc_value[9] = d[509] ^ d[507] ^ d[504] ^ d[502] ^ d[499] ^ d[498] ^ d[494] ^ d[493] ^ d[491] ^ d[488] ^ d[487] ^ d[485] ^ d[482] ^ d[481] ^ d[480] ^ d[479] ^ d[478] ^ d[474] ^ d[471] ^ d[469] ^ d[467] ^ d[466] ^ d[465] ^ d[464] ^ d[463] ^ d[461] ^ d[459] ^ d[456] ^ d[454] ^ d[452] ^ d[451] ^ d[448] ^ d[445] ^ d[442] ^ d[436] ^ d[434] ^ d[433] ^ d[432] ^ d[430] ^ d[427] ^ d[425] ^ d[424] ^ d[423] ^ d[419] ^ d[418] ^ d[416] ^ d[415] ^ d[413] ^ d[411] ^ d[410] ^ d[409] ^ d[404] ^ d[403] ^ d[402] ^ d[401] ^ d[397] ^ d[394] ^ d[391] ^ d[390] ^ d[389] ^ d[388] ^ d[385] ^ d[384] ^ d[382] ^ d[381] ^ d[380] ^ d[379] ^ d[378] ^ d[375] ^ d[374] ^ d[370] ^ d[368] ^ d[367] ^ d[365] ^ d[363] ^ d[362] ^ d[361] ^ d[360] ^ d[358] ^ d[357] ^ d[356] ^ d[355] ^ d[350] ^ d[346] ^ d[338] ^ d[337] ^ d[333] ^ d[330] ^ d[329] ^ d[326] ^ d[324] ^ d[323] ^ d[322] ^ d[319] ^ d[318] ^ d[316] ^ d[315] ^ d[313] ^ d[312] ^ d[309] ^ d[308] ^ d[306] ^ d[305] ^ d[304] ^ d[302] ^ d[300] ^ d[297] ^ d[296] ^ d[295] ^ d[293] ^ d[290] ^ d[287] ^ d[285] ^ d[283] ^ d[282] ^ d[281] ^ d[280] ^ d[278] ^ d[276] ^ d[275] ^ d[274] ^ d[272] ^ d[268] ^ d[266] ^ d[265] ^ d[264] ^ d[263] ^ d[262] ^ d[261] ^ d[260] ^ d[259] ^ d[258] ^ d[257] ^ d[256] ^ d[255] ^ d[254] ^ d[251] ^ d[249] ^ d[248] ^ d[247] ^ d[246] ^ d[243] ^ d[239] ^ d[238] ^ d[236] ^ d[235] ^ d[234] ^ d[233] ^ d[229] ^ d[228] ^ d[227] ^ d[226] ^ d[224] ^ d[222] ^ d[221] ^ d[219] ^ d[217] ^ d[216] ^ d[213] ^ d[211] ^ d[210] ^ d[206] ^ d[203] ^ d[202] ^ d[201] ^ d[200] ^ d[198] ^ d[187] ^ d[186] ^ d[185] ^ d[183] ^ d[181] ^ d[179] ^ d[178] ^ d[177] ^ d[174] ^ d[172] ^ d[171] ^ d[169] ^ d[168] ^ d[167] ^ d[166] ^ d[165] ^ d[164] ^ d[163] ^ d[162] ^ d[161] ^ d[159] ^ d[158] ^ d[157] ^ d[156] ^ d[155] ^ d[154] ^ d[153] ^ d[152] ^ d[151] ^ d[149] ^ d[147] ^ d[143] ^ d[142] ^ d[140] ^ d[138] ^ d[136] ^ d[131] ^ d[129] ^ d[127] ^ d[121] ^ d[120] ^ d[119] ^ d[117] ^ d[115] ^ d[114] ^ d[113] ^ d[110] ^ d[108] ^ d[106] ^ d[104] ^ d[102] ^ d[98] ^ d[96] ^ d[89] ^ d[88] ^ d[86] ^ d[85] ^ d[84] ^ d[83] ^ d[81] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[76] ^ d[74] ^ d[71] ^ d[70] ^ d[69] ^ d[68] ^ d[67] ^ d[66] ^ d[64] ^ d[61] ^ d[60] ^ d[58] ^ d[55] ^ d[53] ^ d[52] ^ d[51] ^ d[47] ^ d[46] ^ d[44] ^ d[43] ^ d[41] ^ d[39] ^ d[38] ^ d[36] ^ d[35] ^ d[34] ^ d[33] ^ d[32] ^ d[29] ^ d[24] ^ d[23] ^ d[18] ^ d[13] ^ d[12] ^ d[11] ^ d[9] ^ d[5] ^ d[4] ^ d[2] ^ d[1] ^ c[0] ^ c[1] ^ c[2] ^ c[5] ^ c[7] ^ c[8] ^ c[11] ^ c[13] ^ c[14] ^ c[18] ^ c[19] ^ c[22] ^ c[24] ^ c[27] ^ c[29];
    stage_2_crc_value[10] = d[511] ^ d[507] ^ d[506] ^ d[505] ^ d[503] ^ d[502] ^ d[501] ^ d[499] ^ d[493] ^ d[491] ^ d[490] ^ d[477] ^ d[476] ^ d[475] ^ d[467] ^ d[466] ^ d[461] ^ d[460] ^ d[458] ^ d[457] ^ d[455] ^ d[453] ^ d[450] ^ d[448] ^ d[446] ^ d[444] ^ d[443] ^ d[436] ^ d[435] ^ d[431] ^ d[428] ^ d[426] ^ d[425] ^ d[422] ^ d[420] ^ d[418] ^ d[417] ^ d[411] ^ d[410] ^ d[409] ^ d[408] ^ d[407] ^ d[403] ^ d[402] ^ d[400] ^ d[399] ^ d[396] ^ d[395] ^ d[393] ^ d[389] ^ d[388] ^ d[387] ^ d[385] ^ d[383] ^ d[382] ^ d[380] ^ d[379] ^ d[378] ^ d[375] ^ d[374] ^ d[372] ^ d[371] ^ d[364] ^ d[361] ^ d[356] ^ d[353] ^ d[351] ^ d[349] ^ d[348] ^ d[345] ^ d[344] ^ d[342] ^ d[341] ^ d[337] ^ d[335] ^ d[333] ^ d[331] ^ d[330] ^ d[328] ^ d[325] ^ d[324] ^ d[323] ^ d[322] ^ d[321] ^ d[318] ^ d[316] ^ d[315] ^ d[314] ^ d[313] ^ d[312] ^ d[307] ^ d[306] ^ d[302] ^ d[301] ^ d[300] ^ d[299] ^ d[295] ^ d[292] ^ d[291] ^ d[290] ^ d[287] ^ d[284] ^ d[282] ^ d[281] ^ d[275] ^ d[274] ^ d[268] ^ d[267] ^ d[266] ^ d[263] ^ d[262] ^ d[260] ^ d[258] ^ d[256] ^ d[250] ^ d[249] ^ d[247] ^ d[244] ^ d[243] ^ d[240] ^ d[239] ^ d[236] ^ d[235] ^ d[229] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[222] ^ d[220] ^ d[218] ^ d[217] ^ d[216] ^ d[211] ^ d[210] ^ d[209] ^ d[208] ^ d[204] ^ d[198] ^ d[197] ^ d[194] ^ d[193] ^ d[192] ^ d[191] ^ d[190] ^ d[187] ^ d[184] ^ d[183] ^ d[180] ^ d[179] ^ d[178] ^ d[175] ^ d[173] ^ d[171] ^ d[168] ^ d[165] ^ d[164] ^ d[163] ^ d[161] ^ d[160] ^ d[159] ^ d[157] ^ d[154] ^ d[153] ^ d[152] ^ d[151] ^ d[150] ^ d[149] ^ d[148] ^ d[141] ^ d[139] ^ d[136] ^ d[135] ^ d[134] ^ d[130] ^ d[127] ^ d[126] ^ d[125] ^ d[123] ^ d[122] ^ d[121] ^ d[120] ^ d[119] ^ d[117] ^ d[115] ^ d[113] ^ d[110] ^ d[109] ^ d[107] ^ d[106] ^ d[105] ^ d[104] ^ d[101] ^ d[98] ^ d[96] ^ d[95] ^ d[94] ^ d[90] ^ d[89] ^ d[86] ^ d[83] ^ d[80] ^ d[78] ^ d[77] ^ d[75] ^ d[73] ^ d[71] ^ d[70] ^ d[69] ^ d[66] ^ d[63] ^ d[62] ^ d[60] ^ d[59] ^ d[58] ^ d[56] ^ d[55] ^ d[52] ^ d[50] ^ d[42] ^ d[40] ^ d[39] ^ d[36] ^ d[35] ^ d[33] ^ d[32] ^ d[31] ^ d[29] ^ d[28] ^ d[26] ^ d[19] ^ d[16] ^ d[14] ^ d[13] ^ d[9] ^ d[5] ^ d[3] ^ d[2] ^ d[0] ^ c[10] ^ c[11] ^ c[13] ^ c[19] ^ c[21] ^ c[22] ^ c[23] ^ c[25] ^ c[26] ^ c[27] ^ c[31];
    stage_2_crc_value[11] = d[511] ^ d[510] ^ d[504] ^ d[503] ^ d[501] ^ d[495] ^ d[493] ^ d[490] ^ d[489] ^ d[488] ^ d[486] ^ d[483] ^ d[482] ^ d[481] ^ d[480] ^ d[479] ^ d[478] ^ d[472] ^ d[470] ^ d[467] ^ d[465] ^ d[464] ^ d[459] ^ d[456] ^ d[454] ^ d[452] ^ d[451] ^ d[450] ^ d[448] ^ d[447] ^ d[445] ^ d[434] ^ d[433] ^ d[432] ^ d[429] ^ d[427] ^ d[426] ^ d[424] ^ d[423] ^ d[422] ^ d[421] ^ d[416] ^ d[414] ^ d[411] ^ d[410] ^ d[407] ^ d[405] ^ d[403] ^ d[401] ^ d[399] ^ d[398] ^ d[397] ^ d[394] ^ d[393] ^ d[392] ^ d[391] ^ d[389] ^ d[387] ^ d[384] ^ d[383] ^ d[380] ^ d[379] ^ d[378] ^ d[375] ^ d[374] ^ d[373] ^ d[369] ^ d[368] ^ d[366] ^ d[365] ^ d[363] ^ d[359] ^ d[358] ^ d[354] ^ d[353] ^ d[352] ^ d[350] ^ d[348] ^ d[347] ^ d[346] ^ d[344] ^ d[343] ^ d[341] ^ d[339] ^ d[337] ^ d[336] ^ d[335] ^ d[333] ^ d[332] ^ d[331] ^ d[329] ^ d[328] ^ d[327] ^ d[326] ^ d[325] ^ d[324] ^ d[323] ^ d[321] ^ d[320] ^ d[318] ^ d[316] ^ d[314] ^ d[313] ^ d[312] ^ d[310] ^ d[309] ^ d[308] ^ d[307] ^ d[305] ^ d[301] ^ d[299] ^ d[298] ^ d[297] ^ d[295] ^ d[294] ^ d[293] ^ d[291] ^ d[290] ^ d[287] ^ d[286] ^ d[285] ^ d[282] ^ d[279] ^ d[277] ^ d[275] ^ d[274] ^ d[273] ^ d[267] ^ d[265] ^ d[263] ^ d[255] ^ d[252] ^ d[251] ^ d[250] ^ d[245] ^ d[244] ^ d[243] ^ d[241] ^ d[240] ^ d[236] ^ d[234] ^ d[228] ^ d[225] ^ d[223] ^ d[221] ^ d[219] ^ d[218] ^ d[217] ^ d[216] ^ d[214] ^ d[211] ^ d[208] ^ d[207] ^ d[205] ^ d[203] ^ d[202] ^ d[201] ^ d[197] ^ d[195] ^ d[190] ^ d[186] ^ d[185] ^ d[184] ^ d[183] ^ d[182] ^ d[181] ^ d[180] ^ d[179] ^ d[176] ^ d[174] ^ d[171] ^ d[170] ^ d[167] ^ d[165] ^ d[164] ^ d[160] ^ d[156] ^ d[154] ^ d[153] ^ d[152] ^ d[150] ^ d[144] ^ d[143] ^ d[142] ^ d[140] ^ d[134] ^ d[132] ^ d[131] ^ d[125] ^ d[124] ^ d[122] ^ d[121] ^ d[120] ^ d[119] ^ d[117] ^ d[113] ^ d[108] ^ d[107] ^ d[105] ^ d[104] ^ d[103] ^ d[102] ^ d[101] ^ d[98] ^ d[94] ^ d[91] ^ d[90] ^ d[85] ^ d[83] ^ d[82] ^ d[78] ^ d[76] ^ d[74] ^ d[73] ^ d[71] ^ d[70] ^ d[68] ^ d[66] ^ d[65] ^ d[64] ^ d[59] ^ d[58] ^ d[57] ^ d[56] ^ d[55] ^ d[54] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[45] ^ d[44] ^ d[43] ^ d[41] ^ d[40] ^ d[36] ^ d[33] ^ d[31] ^ d[28] ^ d[27] ^ d[26] ^ d[25] ^ d[24] ^ d[20] ^ d[17] ^ d[16] ^ d[15] ^ d[14] ^ d[12] ^ d[9] ^ d[4] ^ d[3] ^ d[1] ^ d[0] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[6] ^ c[8] ^ c[9] ^ c[10] ^ c[13] ^ c[15] ^ c[21] ^ c[23] ^ c[24] ^ c[30] ^ c[31];
    stage_2_crc_value[12] = d[510] ^ d[508] ^ d[507] ^ d[506] ^ d[505] ^ d[504] ^ d[501] ^ d[500] ^ d[496] ^ d[495] ^ d[493] ^ d[492] ^ d[488] ^ d[487] ^ d[486] ^ d[484] ^ d[477] ^ d[476] ^ d[473] ^ d[472] ^ d[471] ^ d[470] ^ d[466] ^ d[464] ^ d[462] ^ d[461] ^ d[460] ^ d[458] ^ d[457] ^ d[455] ^ d[453] ^ d[451] ^ d[450] ^ d[446] ^ d[444] ^ d[437] ^ d[436] ^ d[435] ^ d[430] ^ d[428] ^ d[427] ^ d[425] ^ d[423] ^ d[419] ^ d[418] ^ d[417] ^ d[416] ^ d[415] ^ d[414] ^ d[411] ^ d[409] ^ d[407] ^ d[406] ^ d[405] ^ d[402] ^ d[396] ^ d[395] ^ d[394] ^ d[391] ^ d[387] ^ d[386] ^ d[385] ^ d[384] ^ d[380] ^ d[379] ^ d[378] ^ d[375] ^ d[372] ^ d[370] ^ d[368] ^ d[367] ^ d[364] ^ d[363] ^ d[362] ^ d[360] ^ d[358] ^ d[357] ^ d[355] ^ d[354] ^ d[351] ^ d[341] ^ d[340] ^ d[339] ^ d[336] ^ d[335] ^ d[332] ^ d[330] ^ d[329] ^ d[326] ^ d[325] ^ d[324] ^ d[320] ^ d[318] ^ d[314] ^ d[313] ^ d[312] ^ d[311] ^ d[308] ^ d[306] ^ d[305] ^ d[303] ^ d[297] ^ d[291] ^ d[290] ^ d[280] ^ d[279] ^ d[278] ^ d[277] ^ d[275] ^ d[273] ^ d[269] ^ d[266] ^ d[265] ^ d[261] ^ d[259] ^ d[257] ^ d[256] ^ d[255] ^ d[253] ^ d[251] ^ d[248] ^ d[246] ^ d[245] ^ d[244] ^ d[243] ^ d[242] ^ d[241] ^ d[235] ^ d[234] ^ d[230] ^ d[229] ^ d[228] ^ d[227] ^ d[222] ^ d[220] ^ d[219] ^ d[218] ^ d[217] ^ d[216] ^ d[215] ^ d[214] ^ d[210] ^ d[207] ^ d[206] ^ d[204] ^ d[201] ^ d[199] ^ d[197] ^ d[196] ^ d[194] ^ d[193] ^ d[192] ^ d[190] ^ d[188] ^ d[187] ^ d[185] ^ d[184] ^ d[181] ^ d[180] ^ d[177] ^ d[175] ^ d[170] ^ d[169] ^ d[168] ^ d[167] ^ d[165] ^ d[162] ^ d[158] ^ d[157] ^ d[156] ^ d[154] ^ d[153] ^ d[149] ^ d[145] ^ d[141] ^ d[137] ^ d[136] ^ d[134] ^ d[133] ^ d[128] ^ d[127] ^ d[122] ^ d[121] ^ d[120] ^ d[119] ^ d[117] ^ d[116] ^ d[113] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[105] ^ d[102] ^ d[101] ^ d[98] ^ d[97] ^ d[96] ^ d[94] ^ d[92] ^ d[91] ^ d[87] ^ d[86] ^ d[85] ^ d[82] ^ d[81] ^ d[77] ^ d[75] ^ d[74] ^ d[73] ^ d[71] ^ d[69] ^ d[68] ^ d[63] ^ d[61] ^ d[59] ^ d[57] ^ d[56] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[50] ^ d[49] ^ d[47] ^ d[46] ^ d[42] ^ d[41] ^ d[31] ^ d[30] ^ d[27] ^ d[24] ^ d[21] ^ d[18] ^ d[17] ^ d[15] ^ d[13] ^ d[12] ^ d[9] ^ d[6] ^ d[5] ^ d[4] ^ d[2] ^ d[1] ^ d[0] ^ c[4] ^ c[6] ^ c[7] ^ c[8] ^ c[12] ^ c[13] ^ c[15] ^ c[16] ^ c[20] ^ c[21] ^ c[24] ^ c[25] ^ c[26] ^ c[27] ^ c[28] ^ c[30];
    stage_2_crc_value[13] = d[511] ^ d[509] ^ d[508] ^ d[507] ^ d[506] ^ d[505] ^ d[502] ^ d[501] ^ d[497] ^ d[496] ^ d[494] ^ d[493] ^ d[489] ^ d[488] ^ d[487] ^ d[485] ^ d[478] ^ d[477] ^ d[474] ^ d[473] ^ d[472] ^ d[471] ^ d[467] ^ d[465] ^ d[463] ^ d[462] ^ d[461] ^ d[459] ^ d[458] ^ d[456] ^ d[454] ^ d[452] ^ d[451] ^ d[447] ^ d[445] ^ d[438] ^ d[437] ^ d[436] ^ d[431] ^ d[429] ^ d[428] ^ d[426] ^ d[424] ^ d[420] ^ d[419] ^ d[418] ^ d[417] ^ d[416] ^ d[415] ^ d[412] ^ d[410] ^ d[408] ^ d[407] ^ d[406] ^ d[403] ^ d[397] ^ d[396] ^ d[395] ^ d[392] ^ d[388] ^ d[387] ^ d[386] ^ d[385] ^ d[381] ^ d[380] ^ d[379] ^ d[376] ^ d[373] ^ d[371] ^ d[369] ^ d[368] ^ d[365] ^ d[364] ^ d[363] ^ d[361] ^ d[359] ^ d[358] ^ d[356] ^ d[355] ^ d[352] ^ d[342] ^ d[341] ^ d[340] ^ d[337] ^ d[336] ^ d[333] ^ d[331] ^ d[330] ^ d[327] ^ d[326] ^ d[325] ^ d[321] ^ d[319] ^ d[315] ^ d[314] ^ d[313] ^ d[312] ^ d[309] ^ d[307] ^ d[306] ^ d[304] ^ d[298] ^ d[292] ^ d[291] ^ d[281] ^ d[280] ^ d[279] ^ d[278] ^ d[276] ^ d[274] ^ d[270] ^ d[267] ^ d[266] ^ d[262] ^ d[260] ^ d[258] ^ d[257] ^ d[256] ^ d[254] ^ d[252] ^ d[249] ^ d[247] ^ d[246] ^ d[245] ^ d[244] ^ d[243] ^ d[242] ^ d[236] ^ d[235] ^ d[231] ^ d[230] ^ d[229] ^ d[228] ^ d[223] ^ d[221] ^ d[220] ^ d[219] ^ d[218] ^ d[217] ^ d[216] ^ d[215] ^ d[211] ^ d[208] ^ d[207] ^ d[205] ^ d[202] ^ d[200] ^ d[198] ^ d[197] ^ d[195] ^ d[194] ^ d[193] ^ d[191] ^ d[189] ^ d[188] ^ d[186] ^ d[185] ^ d[182] ^ d[181] ^ d[178] ^ d[176] ^ d[171] ^ d[170] ^ d[169] ^ d[168] ^ d[166] ^ d[163] ^ d[159] ^ d[158] ^ d[157] ^ d[155] ^ d[154] ^ d[150] ^ d[146] ^ d[142] ^ d[138] ^ d[137] ^ d[135] ^ d[134] ^ d[129] ^ d[128] ^ d[123] ^ d[122] ^ d[121] ^ d[120] ^ d[118] ^ d[117] ^ d[114] ^ d[112] ^ d[111] ^ d[110] ^ d[109] ^ d[106] ^ d[103] ^ d[102] ^ d[99] ^ d[98] ^ d[97] ^ d[95] ^ d[93] ^ d[92] ^ d[88] ^ d[87] ^ d[86] ^ d[83] ^ d[82] ^ d[78] ^ d[76] ^ d[75] ^ d[74] ^ d[72] ^ d[70] ^ d[69] ^ d[64] ^ d[62] ^ d[60] ^ d[58] ^ d[57] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[43] ^ d[42] ^ d[32] ^ d[31] ^ d[28] ^ d[25] ^ d[22] ^ d[19] ^ d[18] ^ d[16] ^ d[14] ^ d[13] ^ d[10] ^ d[7] ^ d[6] ^ d[5] ^ d[3] ^ d[2] ^ d[1] ^ c[5] ^ c[7] ^ c[8] ^ c[9] ^ c[13] ^ c[14] ^ c[16] ^ c[17] ^ c[21] ^ c[22] ^ c[25] ^ c[26] ^ c[27] ^ c[28] ^ c[29] ^ c[31];
    stage_2_crc_value[14] = d[510] ^ d[509] ^ d[508] ^ d[507] ^ d[506] ^ d[503] ^ d[502] ^ d[498] ^ d[497] ^ d[495] ^ d[494] ^ d[490] ^ d[489] ^ d[488] ^ d[486] ^ d[479] ^ d[478] ^ d[475] ^ d[474] ^ d[473] ^ d[472] ^ d[468] ^ d[466] ^ d[464] ^ d[463] ^ d[462] ^ d[460] ^ d[459] ^ d[457] ^ d[455] ^ d[453] ^ d[452] ^ d[448] ^ d[446] ^ d[439] ^ d[438] ^ d[437] ^ d[432] ^ d[430] ^ d[429] ^ d[427] ^ d[425] ^ d[421] ^ d[420] ^ d[419] ^ d[418] ^ d[417] ^ d[416] ^ d[413] ^ d[411] ^ d[409] ^ d[408] ^ d[407] ^ d[404] ^ d[398] ^ d[397] ^ d[396] ^ d[393] ^ d[389] ^ d[388] ^ d[387] ^ d[386] ^ d[382] ^ d[381] ^ d[380] ^ d[377] ^ d[374] ^ d[372] ^ d[370] ^ d[369] ^ d[366] ^ d[365] ^ d[364] ^ d[362] ^ d[360] ^ d[359] ^ d[357] ^ d[356] ^ d[353] ^ d[343] ^ d[342] ^ d[341] ^ d[338] ^ d[337] ^ d[334] ^ d[332] ^ d[331] ^ d[328] ^ d[327] ^ d[326] ^ d[322] ^ d[320] ^ d[316] ^ d[315] ^ d[314] ^ d[313] ^ d[310] ^ d[308] ^ d[307] ^ d[305] ^ d[299] ^ d[293] ^ d[292] ^ d[282] ^ d[281] ^ d[280] ^ d[279] ^ d[277] ^ d[275] ^ d[271] ^ d[268] ^ d[267] ^ d[263] ^ d[261] ^ d[259] ^ d[258] ^ d[257] ^ d[255] ^ d[253] ^ d[250] ^ d[248] ^ d[247] ^ d[246] ^ d[245] ^ d[244] ^ d[243] ^ d[237] ^ d[236] ^ d[232] ^ d[231] ^ d[230] ^ d[229] ^ d[224] ^ d[222] ^ d[221] ^ d[220] ^ d[219] ^ d[218] ^ d[217] ^ d[216] ^ d[212] ^ d[209] ^ d[208] ^ d[206] ^ d[203] ^ d[201] ^ d[199] ^ d[198] ^ d[196] ^ d[195] ^ d[194] ^ d[192] ^ d[190] ^ d[189] ^ d[187] ^ d[186] ^ d[183] ^ d[182] ^ d[179] ^ d[177] ^ d[172] ^ d[171] ^ d[170] ^ d[169] ^ d[167] ^ d[164] ^ d[160] ^ d[159] ^ d[158] ^ d[156] ^ d[155] ^ d[151] ^ d[147] ^ d[143] ^ d[139] ^ d[138] ^ d[136] ^ d[135] ^ d[130] ^ d[129] ^ d[124] ^ d[123] ^ d[122] ^ d[121] ^ d[119] ^ d[118] ^ d[115] ^ d[113] ^ d[112] ^ d[111] ^ d[110] ^ d[107] ^ d[104] ^ d[103] ^ d[100] ^ d[99] ^ d[98] ^ d[96] ^ d[94] ^ d[93] ^ d[89] ^ d[88] ^ d[87] ^ d[84] ^ d[83] ^ d[79] ^ d[77] ^ d[76] ^ d[75] ^ d[73] ^ d[71] ^ d[70] ^ d[65] ^ d[63] ^ d[61] ^ d[59] ^ d[58] ^ d[56] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[49] ^ d[48] ^ d[44] ^ d[43] ^ d[33] ^ d[32] ^ d[29] ^ d[26] ^ d[23] ^ d[20] ^ d[19] ^ d[17] ^ d[15] ^ d[14] ^ d[11] ^ d[8] ^ d[7] ^ d[6] ^ d[4] ^ d[3] ^ d[2] ^ c[6] ^ c[8] ^ c[9] ^ c[10] ^ c[14] ^ c[15] ^ c[17] ^ c[18] ^ c[22] ^ c[23] ^ c[26] ^ c[27] ^ c[28] ^ c[29] ^ c[30];
    stage_2_crc_value[15] = d[511] ^ d[510] ^ d[509] ^ d[508] ^ d[507] ^ d[504] ^ d[503] ^ d[499] ^ d[498] ^ d[496] ^ d[495] ^ d[491] ^ d[490] ^ d[489] ^ d[487] ^ d[480] ^ d[479] ^ d[476] ^ d[475] ^ d[474] ^ d[473] ^ d[469] ^ d[467] ^ d[465] ^ d[464] ^ d[463] ^ d[461] ^ d[460] ^ d[458] ^ d[456] ^ d[454] ^ d[453] ^ d[449] ^ d[447] ^ d[440] ^ d[439] ^ d[438] ^ d[433] ^ d[431] ^ d[430] ^ d[428] ^ d[426] ^ d[422] ^ d[421] ^ d[420] ^ d[419] ^ d[418] ^ d[417] ^ d[414] ^ d[412] ^ d[410] ^ d[409] ^ d[408] ^ d[405] ^ d[399] ^ d[398] ^ d[397] ^ d[394] ^ d[390] ^ d[389] ^ d[388] ^ d[387] ^ d[383] ^ d[382] ^ d[381] ^ d[378] ^ d[375] ^ d[373] ^ d[371] ^ d[370] ^ d[367] ^ d[366] ^ d[365] ^ d[363] ^ d[361] ^ d[360] ^ d[358] ^ d[357] ^ d[354] ^ d[344] ^ d[343] ^ d[342] ^ d[339] ^ d[338] ^ d[335] ^ d[333] ^ d[332] ^ d[329] ^ d[328] ^ d[327] ^ d[323] ^ d[321] ^ d[317] ^ d[316] ^ d[315] ^ d[314] ^ d[311] ^ d[309] ^ d[308] ^ d[306] ^ d[300] ^ d[294] ^ d[293] ^ d[283] ^ d[282] ^ d[281] ^ d[280] ^ d[278] ^ d[276] ^ d[272] ^ d[269] ^ d[268] ^ d[264] ^ d[262] ^ d[260] ^ d[259] ^ d[258] ^ d[256] ^ d[254] ^ d[251] ^ d[249] ^ d[248] ^ d[247] ^ d[246] ^ d[245] ^ d[244] ^ d[238] ^ d[237] ^ d[233] ^ d[232] ^ d[231] ^ d[230] ^ d[225] ^ d[223] ^ d[222] ^ d[221] ^ d[220] ^ d[219] ^ d[218] ^ d[217] ^ d[213] ^ d[210] ^ d[209] ^ d[207] ^ d[204] ^ d[202] ^ d[200] ^ d[199] ^ d[197] ^ d[196] ^ d[195] ^ d[193] ^ d[191] ^ d[190] ^ d[188] ^ d[187] ^ d[184] ^ d[183] ^ d[180] ^ d[178] ^ d[173] ^ d[172] ^ d[171] ^ d[170] ^ d[168] ^ d[165] ^ d[161] ^ d[160] ^ d[159] ^ d[157] ^ d[156] ^ d[152] ^ d[148] ^ d[144] ^ d[140] ^ d[139] ^ d[137] ^ d[136] ^ d[131] ^ d[130] ^ d[125] ^ d[124] ^ d[123] ^ d[122] ^ d[120] ^ d[119] ^ d[116] ^ d[114] ^ d[113] ^ d[112] ^ d[111] ^ d[108] ^ d[105] ^ d[104] ^ d[101] ^ d[100] ^ d[99] ^ d[97] ^ d[95] ^ d[94] ^ d[90] ^ d[89] ^ d[88] ^ d[85] ^ d[84] ^ d[80] ^ d[78] ^ d[77] ^ d[76] ^ d[74] ^ d[72] ^ d[71] ^ d[66] ^ d[64] ^ d[62] ^ d[60] ^ d[59] ^ d[57] ^ d[56] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[50] ^ d[49] ^ d[45] ^ d[44] ^ d[34] ^ d[33] ^ d[30] ^ d[27] ^ d[24] ^ d[21] ^ d[20] ^ d[18] ^ d[16] ^ d[15] ^ d[12] ^ d[9] ^ d[8] ^ d[7] ^ d[5] ^ d[4] ^ d[3] ^ c[0] ^ c[7] ^ c[9] ^ c[10] ^ c[11] ^ c[15] ^ c[16] ^ c[18] ^ c[19] ^ c[23] ^ c[24] ^ c[27] ^ c[28] ^ c[29] ^ c[30] ^ c[31];
    stage_2_crc_value[16] = d[509] ^ d[507] ^ d[506] ^ d[505] ^ d[504] ^ d[502] ^ d[501] ^ d[499] ^ d[497] ^ d[496] ^ d[495] ^ d[494] ^ d[493] ^ d[489] ^ d[486] ^ d[483] ^ d[482] ^ d[479] ^ d[475] ^ d[474] ^ d[472] ^ d[466] ^ d[459] ^ d[458] ^ d[457] ^ d[455] ^ d[454] ^ d[452] ^ d[449] ^ d[444] ^ d[441] ^ d[440] ^ d[439] ^ d[437] ^ d[436] ^ d[433] ^ d[432] ^ d[431] ^ d[429] ^ d[427] ^ d[424] ^ d[423] ^ d[421] ^ d[420] ^ d[416] ^ d[415] ^ d[414] ^ d[413] ^ d[412] ^ d[411] ^ d[410] ^ d[408] ^ d[407] ^ d[406] ^ d[405] ^ d[404] ^ d[396] ^ d[395] ^ d[393] ^ d[392] ^ d[389] ^ d[387] ^ d[386] ^ d[384] ^ d[383] ^ d[382] ^ d[381] ^ d[379] ^ d[378] ^ d[371] ^ d[369] ^ d[367] ^ d[364] ^ d[363] ^ d[361] ^ d[357] ^ d[355] ^ d[353] ^ d[349] ^ d[348] ^ d[347] ^ d[343] ^ d[342] ^ d[341] ^ d[340] ^ d[338] ^ d[337] ^ d[336] ^ d[335] ^ d[330] ^ d[329] ^ d[327] ^ d[324] ^ d[321] ^ d[320] ^ d[319] ^ d[316] ^ d[307] ^ d[305] ^ d[303] ^ d[302] ^ d[301] ^ d[300] ^ d[299] ^ d[298] ^ d[297] ^ d[296] ^ d[292] ^ d[290] ^ d[288] ^ d[287] ^ d[286] ^ d[284] ^ d[282] ^ d[281] ^ d[276] ^ d[274] ^ d[270] ^ d[268] ^ d[264] ^ d[263] ^ d[260] ^ d[250] ^ d[249] ^ d[247] ^ d[246] ^ d[245] ^ d[243] ^ d[239] ^ d[238] ^ d[237] ^ d[233] ^ d[232] ^ d[231] ^ d[230] ^ d[228] ^ d[227] ^ d[223] ^ d[222] ^ d[221] ^ d[220] ^ d[219] ^ d[218] ^ d[216] ^ d[212] ^ d[211] ^ d[209] ^ d[207] ^ d[205] ^ d[202] ^ d[200] ^ d[199] ^ d[196] ^ d[193] ^ d[190] ^ d[189] ^ d[186] ^ d[185] ^ d[184] ^ d[183] ^ d[182] ^ d[181] ^ d[179] ^ d[174] ^ d[173] ^ d[170] ^ d[167] ^ d[160] ^ d[157] ^ d[156] ^ d[155] ^ d[153] ^ d[151] ^ d[145] ^ d[144] ^ d[143] ^ d[141] ^ d[140] ^ d[138] ^ d[136] ^ d[135] ^ d[134] ^ d[131] ^ d[128] ^ d[127] ^ d[124] ^ d[121] ^ d[120] ^ d[119] ^ d[118] ^ d[116] ^ d[115] ^ d[112] ^ d[111] ^ d[110] ^ d[109] ^ d[105] ^ d[104] ^ d[103] ^ d[102] ^ d[100] ^ d[99] ^ d[97] ^ d[94] ^ d[91] ^ d[90] ^ d[89] ^ d[87] ^ d[86] ^ d[84] ^ d[83] ^ d[82] ^ d[78] ^ d[77] ^ d[75] ^ d[68] ^ d[66] ^ d[57] ^ d[56] ^ d[51] ^ d[48] ^ d[47] ^ d[46] ^ d[44] ^ d[37] ^ d[35] ^ d[32] ^ d[30] ^ d[29] ^ d[26] ^ d[24] ^ d[22] ^ d[21] ^ d[19] ^ d[17] ^ d[13] ^ d[12] ^ d[8] ^ d[5] ^ d[4] ^ d[0] ^ c[2] ^ c[3] ^ c[6] ^ c[9] ^ c[13] ^ c[14] ^ c[15] ^ c[16] ^ c[17] ^ c[19] ^ c[21] ^ c[22] ^ c[24] ^ c[25] ^ c[26] ^ c[27] ^ c[29];
    stage_2_crc_value[17] = d[510] ^ d[508] ^ d[507] ^ d[506] ^ d[505] ^ d[503] ^ d[502] ^ d[500] ^ d[498] ^ d[497] ^ d[496] ^ d[495] ^ d[494] ^ d[490] ^ d[487] ^ d[484] ^ d[483] ^ d[480] ^ d[476] ^ d[475] ^ d[473] ^ d[467] ^ d[460] ^ d[459] ^ d[458] ^ d[456] ^ d[455] ^ d[453] ^ d[450] ^ d[445] ^ d[442] ^ d[441] ^ d[440] ^ d[438] ^ d[437] ^ d[434] ^ d[433] ^ d[432] ^ d[430] ^ d[428] ^ d[425] ^ d[424] ^ d[422] ^ d[421] ^ d[417] ^ d[416] ^ d[415] ^ d[414] ^ d[413] ^ d[412] ^ d[411] ^ d[409] ^ d[408] ^ d[407] ^ d[406] ^ d[405] ^ d[397] ^ d[396] ^ d[394] ^ d[393] ^ d[390] ^ d[388] ^ d[387] ^ d[385] ^ d[384] ^ d[383] ^ d[382] ^ d[380] ^ d[379] ^ d[372] ^ d[370] ^ d[368] ^ d[365] ^ d[364] ^ d[362] ^ d[358] ^ d[356] ^ d[354] ^ d[350] ^ d[349] ^ d[348] ^ d[344] ^ d[343] ^ d[342] ^ d[341] ^ d[339] ^ d[338] ^ d[337] ^ d[336] ^ d[331] ^ d[330] ^ d[328] ^ d[325] ^ d[322] ^ d[321] ^ d[320] ^ d[317] ^ d[308] ^ d[306] ^ d[304] ^ d[303] ^ d[302] ^ d[301] ^ d[300] ^ d[299] ^ d[298] ^ d[297] ^ d[293] ^ d[291] ^ d[289] ^ d[288] ^ d[287] ^ d[285] ^ d[283] ^ d[282] ^ d[277] ^ d[275] ^ d[271] ^ d[269] ^ d[265] ^ d[264] ^ d[261] ^ d[251] ^ d[250] ^ d[248] ^ d[247] ^ d[246] ^ d[244] ^ d[240] ^ d[239] ^ d[238] ^ d[234] ^ d[233] ^ d[232] ^ d[231] ^ d[229] ^ d[228] ^ d[224] ^ d[223] ^ d[222] ^ d[221] ^ d[220] ^ d[219] ^ d[217] ^ d[213] ^ d[212] ^ d[210] ^ d[208] ^ d[206] ^ d[203] ^ d[201] ^ d[200] ^ d[197] ^ d[194] ^ d[191] ^ d[190] ^ d[187] ^ d[186] ^ d[185] ^ d[184] ^ d[183] ^ d[182] ^ d[180] ^ d[175] ^ d[174] ^ d[171] ^ d[168] ^ d[161] ^ d[158] ^ d[157] ^ d[156] ^ d[154] ^ d[152] ^ d[146] ^ d[145] ^ d[144] ^ d[142] ^ d[141] ^ d[139] ^ d[137] ^ d[136] ^ d[135] ^ d[132] ^ d[129] ^ d[128] ^ d[125] ^ d[122] ^ d[121] ^ d[120] ^ d[119] ^ d[117] ^ d[116] ^ d[113] ^ d[112] ^ d[111] ^ d[110] ^ d[106] ^ d[105] ^ d[104] ^ d[103] ^ d[101] ^ d[100] ^ d[98] ^ d[95] ^ d[92] ^ d[91] ^ d[90] ^ d[88] ^ d[87] ^ d[85] ^ d[84] ^ d[83] ^ d[79] ^ d[78] ^ d[76] ^ d[69] ^ d[67] ^ d[58] ^ d[57] ^ d[52] ^ d[49] ^ d[48] ^ d[47] ^ d[45] ^ d[38] ^ d[36] ^ d[33] ^ d[31] ^ d[30] ^ d[27] ^ d[25] ^ d[23] ^ d[22] ^ d[20] ^ d[18] ^ d[14] ^ d[13] ^ d[9] ^ d[6] ^ d[5] ^ d[1] ^ c[0] ^ c[3] ^ c[4] ^ c[7] ^ c[10] ^ c[14] ^ c[15] ^ c[16] ^ c[17] ^ c[18] ^ c[20] ^ c[22] ^ c[23] ^ c[25] ^ c[26] ^ c[27] ^ c[28] ^ c[30];
    stage_2_crc_value[18] = d[511] ^ d[509] ^ d[508] ^ d[507] ^ d[506] ^ d[504] ^ d[503] ^ d[501] ^ d[499] ^ d[498] ^ d[497] ^ d[496] ^ d[495] ^ d[491] ^ d[488] ^ d[485] ^ d[484] ^ d[481] ^ d[477] ^ d[476] ^ d[474] ^ d[468] ^ d[461] ^ d[460] ^ d[459] ^ d[457] ^ d[456] ^ d[454] ^ d[451] ^ d[446] ^ d[443] ^ d[442] ^ d[441] ^ d[439] ^ d[438] ^ d[435] ^ d[434] ^ d[433] ^ d[431] ^ d[429] ^ d[426] ^ d[425] ^ d[423] ^ d[422] ^ d[418] ^ d[417] ^ d[416] ^ d[415] ^ d[414] ^ d[413] ^ d[412] ^ d[410] ^ d[409] ^ d[408] ^ d[407] ^ d[406] ^ d[398] ^ d[397] ^ d[395] ^ d[394] ^ d[391] ^ d[389] ^ d[388] ^ d[386] ^ d[385] ^ d[384] ^ d[383] ^ d[381] ^ d[380] ^ d[373] ^ d[371] ^ d[369] ^ d[366] ^ d[365] ^ d[363] ^ d[359] ^ d[357] ^ d[355] ^ d[351] ^ d[350] ^ d[349] ^ d[345] ^ d[344] ^ d[343] ^ d[342] ^ d[340] ^ d[339] ^ d[338] ^ d[337] ^ d[332] ^ d[331] ^ d[329] ^ d[326] ^ d[323] ^ d[322] ^ d[321] ^ d[318] ^ d[309] ^ d[307] ^ d[305] ^ d[304] ^ d[303] ^ d[302] ^ d[301] ^ d[300] ^ d[299] ^ d[298] ^ d[294] ^ d[292] ^ d[290] ^ d[289] ^ d[288] ^ d[286] ^ d[284] ^ d[283] ^ d[278] ^ d[276] ^ d[272] ^ d[270] ^ d[266] ^ d[265] ^ d[262] ^ d[252] ^ d[251] ^ d[249] ^ d[248] ^ d[247] ^ d[245] ^ d[241] ^ d[240] ^ d[239] ^ d[235] ^ d[234] ^ d[233] ^ d[232] ^ d[230] ^ d[229] ^ d[225] ^ d[224] ^ d[223] ^ d[222] ^ d[221] ^ d[220] ^ d[218] ^ d[214] ^ d[213] ^ d[211] ^ d[209] ^ d[207] ^ d[204] ^ d[202] ^ d[201] ^ d[198] ^ d[195] ^ d[192] ^ d[191] ^ d[188] ^ d[187] ^ d[186] ^ d[185] ^ d[184] ^ d[183] ^ d[181] ^ d[176] ^ d[175] ^ d[172] ^ d[169] ^ d[162] ^ d[159] ^ d[158] ^ d[157] ^ d[155] ^ d[153] ^ d[147] ^ d[146] ^ d[145] ^ d[143] ^ d[142] ^ d[140] ^ d[138] ^ d[137] ^ d[136] ^ d[133] ^ d[130] ^ d[129] ^ d[126] ^ d[123] ^ d[122] ^ d[121] ^ d[120] ^ d[118] ^ d[117] ^ d[114] ^ d[113] ^ d[112] ^ d[111] ^ d[107] ^ d[106] ^ d[105] ^ d[104] ^ d[102] ^ d[101] ^ d[99] ^ d[96] ^ d[93] ^ d[92] ^ d[91] ^ d[89] ^ d[88] ^ d[86] ^ d[85] ^ d[84] ^ d[80] ^ d[79] ^ d[77] ^ d[70] ^ d[68] ^ d[59] ^ d[58] ^ d[53] ^ d[50] ^ d[49] ^ d[48] ^ d[46] ^ d[39] ^ d[37] ^ d[34] ^ d[32] ^ d[31] ^ d[28] ^ d[26] ^ d[24] ^ d[23] ^ d[21] ^ d[19] ^ d[15] ^ d[14] ^ d[10] ^ d[7] ^ d[6] ^ d[2] ^ c[1] ^ c[4] ^ c[5] ^ c[8] ^ c[11] ^ c[15] ^ c[16] ^ c[17] ^ c[18] ^ c[19] ^ c[21] ^ c[23] ^ c[24] ^ c[26] ^ c[27] ^ c[28] ^ c[29] ^ c[31];
    stage_2_crc_value[19] = d[510] ^ d[509] ^ d[508] ^ d[507] ^ d[505] ^ d[504] ^ d[502] ^ d[500] ^ d[499] ^ d[498] ^ d[497] ^ d[496] ^ d[492] ^ d[489] ^ d[486] ^ d[485] ^ d[482] ^ d[478] ^ d[477] ^ d[475] ^ d[469] ^ d[462] ^ d[461] ^ d[460] ^ d[458] ^ d[457] ^ d[455] ^ d[452] ^ d[447] ^ d[444] ^ d[443] ^ d[442] ^ d[440] ^ d[439] ^ d[436] ^ d[435] ^ d[434] ^ d[432] ^ d[430] ^ d[427] ^ d[426] ^ d[424] ^ d[423] ^ d[419] ^ d[418] ^ d[417] ^ d[416] ^ d[415] ^ d[414] ^ d[413] ^ d[411] ^ d[410] ^ d[409] ^ d[408] ^ d[407] ^ d[399] ^ d[398] ^ d[396] ^ d[395] ^ d[392] ^ d[390] ^ d[389] ^ d[387] ^ d[386] ^ d[385] ^ d[384] ^ d[382] ^ d[381] ^ d[374] ^ d[372] ^ d[370] ^ d[367] ^ d[366] ^ d[364] ^ d[360] ^ d[358] ^ d[356] ^ d[352] ^ d[351] ^ d[350] ^ d[346] ^ d[345] ^ d[344] ^ d[343] ^ d[341] ^ d[340] ^ d[339] ^ d[338] ^ d[333] ^ d[332] ^ d[330] ^ d[327] ^ d[324] ^ d[323] ^ d[322] ^ d[319] ^ d[310] ^ d[308] ^ d[306] ^ d[305] ^ d[304] ^ d[303] ^ d[302] ^ d[301] ^ d[300] ^ d[299] ^ d[295] ^ d[293] ^ d[291] ^ d[290] ^ d[289] ^ d[287] ^ d[285] ^ d[284] ^ d[279] ^ d[277] ^ d[273] ^ d[271] ^ d[267] ^ d[266] ^ d[263] ^ d[253] ^ d[252] ^ d[250] ^ d[249] ^ d[248] ^ d[246] ^ d[242] ^ d[241] ^ d[240] ^ d[236] ^ d[235] ^ d[234] ^ d[233] ^ d[231] ^ d[230] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[222] ^ d[221] ^ d[219] ^ d[215] ^ d[214] ^ d[212] ^ d[210] ^ d[208] ^ d[205] ^ d[203] ^ d[202] ^ d[199] ^ d[196] ^ d[193] ^ d[192] ^ d[189] ^ d[188] ^ d[187] ^ d[186] ^ d[185] ^ d[184] ^ d[182] ^ d[177] ^ d[176] ^ d[173] ^ d[170] ^ d[163] ^ d[160] ^ d[159] ^ d[158] ^ d[156] ^ d[154] ^ d[148] ^ d[147] ^ d[146] ^ d[144] ^ d[143] ^ d[141] ^ d[139] ^ d[138] ^ d[137] ^ d[134] ^ d[131] ^ d[130] ^ d[127] ^ d[124] ^ d[123] ^ d[122] ^ d[121] ^ d[119] ^ d[118] ^ d[115] ^ d[114] ^ d[113] ^ d[112] ^ d[108] ^ d[107] ^ d[106] ^ d[105] ^ d[103] ^ d[102] ^ d[100] ^ d[97] ^ d[94] ^ d[93] ^ d[92] ^ d[90] ^ d[89] ^ d[87] ^ d[86] ^ d[85] ^ d[81] ^ d[80] ^ d[78] ^ d[71] ^ d[69] ^ d[60] ^ d[59] ^ d[54] ^ d[51] ^ d[50] ^ d[49] ^ d[47] ^ d[40] ^ d[38] ^ d[35] ^ d[33] ^ d[32] ^ d[29] ^ d[27] ^ d[25] ^ d[24] ^ d[22] ^ d[20] ^ d[16] ^ d[15] ^ d[11] ^ d[8] ^ d[7] ^ d[3] ^ c[2] ^ c[5] ^ c[6] ^ c[9] ^ c[12] ^ c[16] ^ c[17] ^ c[18] ^ c[19] ^ c[20] ^ c[22] ^ c[24] ^ c[25] ^ c[27] ^ c[28] ^ c[29] ^ c[30];
    stage_2_crc_value[20] = d[511] ^ d[510] ^ d[509] ^ d[508] ^ d[506] ^ d[505] ^ d[503] ^ d[501] ^ d[500] ^ d[499] ^ d[498] ^ d[497] ^ d[493] ^ d[490] ^ d[487] ^ d[486] ^ d[483] ^ d[479] ^ d[478] ^ d[476] ^ d[470] ^ d[463] ^ d[462] ^ d[461] ^ d[459] ^ d[458] ^ d[456] ^ d[453] ^ d[448] ^ d[445] ^ d[444] ^ d[443] ^ d[441] ^ d[440] ^ d[437] ^ d[436] ^ d[435] ^ d[433] ^ d[431] ^ d[428] ^ d[427] ^ d[425] ^ d[424] ^ d[420] ^ d[419] ^ d[418] ^ d[417] ^ d[416] ^ d[415] ^ d[414] ^ d[412] ^ d[411] ^ d[410] ^ d[409] ^ d[408] ^ d[400] ^ d[399] ^ d[397] ^ d[396] ^ d[393] ^ d[391] ^ d[390] ^ d[388] ^ d[387] ^ d[386] ^ d[385] ^ d[383] ^ d[382] ^ d[375] ^ d[373] ^ d[371] ^ d[368] ^ d[367] ^ d[365] ^ d[361] ^ d[359] ^ d[357] ^ d[353] ^ d[352] ^ d[351] ^ d[347] ^ d[346] ^ d[345] ^ d[344] ^ d[342] ^ d[341] ^ d[340] ^ d[339] ^ d[334] ^ d[333] ^ d[331] ^ d[328] ^ d[325] ^ d[324] ^ d[323] ^ d[320] ^ d[311] ^ d[309] ^ d[307] ^ d[306] ^ d[305] ^ d[304] ^ d[303] ^ d[302] ^ d[301] ^ d[300] ^ d[296] ^ d[294] ^ d[292] ^ d[291] ^ d[290] ^ d[288] ^ d[286] ^ d[285] ^ d[280] ^ d[278] ^ d[274] ^ d[272] ^ d[268] ^ d[267] ^ d[264] ^ d[254] ^ d[253] ^ d[251] ^ d[250] ^ d[249] ^ d[247] ^ d[243] ^ d[242] ^ d[241] ^ d[237] ^ d[236] ^ d[235] ^ d[234] ^ d[232] ^ d[231] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[222] ^ d[220] ^ d[216] ^ d[215] ^ d[213] ^ d[211] ^ d[209] ^ d[206] ^ d[204] ^ d[203] ^ d[200] ^ d[197] ^ d[194] ^ d[193] ^ d[190] ^ d[189] ^ d[188] ^ d[187] ^ d[186] ^ d[185] ^ d[183] ^ d[178] ^ d[177] ^ d[174] ^ d[171] ^ d[164] ^ d[161] ^ d[160] ^ d[159] ^ d[157] ^ d[155] ^ d[149] ^ d[148] ^ d[147] ^ d[145] ^ d[144] ^ d[142] ^ d[140] ^ d[139] ^ d[138] ^ d[135] ^ d[132] ^ d[131] ^ d[128] ^ d[125] ^ d[124] ^ d[123] ^ d[122] ^ d[120] ^ d[119] ^ d[116] ^ d[115] ^ d[114] ^ d[113] ^ d[109] ^ d[108] ^ d[107] ^ d[106] ^ d[104] ^ d[103] ^ d[101] ^ d[98] ^ d[95] ^ d[94] ^ d[93] ^ d[91] ^ d[90] ^ d[88] ^ d[87] ^ d[86] ^ d[82] ^ d[81] ^ d[79] ^ d[72] ^ d[70] ^ d[61] ^ d[60] ^ d[55] ^ d[52] ^ d[51] ^ d[50] ^ d[48] ^ d[41] ^ d[39] ^ d[36] ^ d[34] ^ d[33] ^ d[30] ^ d[28] ^ d[26] ^ d[25] ^ d[23] ^ d[21] ^ d[17] ^ d[16] ^ d[12] ^ d[9] ^ d[8] ^ d[4] ^ c[3] ^ c[6] ^ c[7] ^ c[10] ^ c[13] ^ c[17] ^ c[18] ^ c[19] ^ c[20] ^ c[21] ^ c[23] ^ c[25] ^ c[26] ^ c[28] ^ c[29] ^ c[30] ^ c[31];
    stage_2_crc_value[21] = d[511] ^ d[510] ^ d[509] ^ d[507] ^ d[506] ^ d[504] ^ d[502] ^ d[501] ^ d[500] ^ d[499] ^ d[498] ^ d[494] ^ d[491] ^ d[488] ^ d[487] ^ d[484] ^ d[480] ^ d[479] ^ d[477] ^ d[471] ^ d[464] ^ d[463] ^ d[462] ^ d[460] ^ d[459] ^ d[457] ^ d[454] ^ d[449] ^ d[446] ^ d[445] ^ d[444] ^ d[442] ^ d[441] ^ d[438] ^ d[437] ^ d[436] ^ d[434] ^ d[432] ^ d[429] ^ d[428] ^ d[426] ^ d[425] ^ d[421] ^ d[420] ^ d[419] ^ d[418] ^ d[417] ^ d[416] ^ d[415] ^ d[413] ^ d[412] ^ d[411] ^ d[410] ^ d[409] ^ d[401] ^ d[400] ^ d[398] ^ d[397] ^ d[394] ^ d[392] ^ d[391] ^ d[389] ^ d[388] ^ d[387] ^ d[386] ^ d[384] ^ d[383] ^ d[376] ^ d[374] ^ d[372] ^ d[369] ^ d[368] ^ d[366] ^ d[362] ^ d[360] ^ d[358] ^ d[354] ^ d[353] ^ d[352] ^ d[348] ^ d[347] ^ d[346] ^ d[345] ^ d[343] ^ d[342] ^ d[341] ^ d[340] ^ d[335] ^ d[334] ^ d[332] ^ d[329] ^ d[326] ^ d[325] ^ d[324] ^ d[321] ^ d[312] ^ d[310] ^ d[308] ^ d[307] ^ d[306] ^ d[305] ^ d[304] ^ d[303] ^ d[302] ^ d[301] ^ d[297] ^ d[295] ^ d[293] ^ d[292] ^ d[291] ^ d[289] ^ d[287] ^ d[286] ^ d[281] ^ d[279] ^ d[275] ^ d[273] ^ d[269] ^ d[268] ^ d[265] ^ d[255] ^ d[254] ^ d[252] ^ d[251] ^ d[250] ^ d[248] ^ d[244] ^ d[243] ^ d[242] ^ d[238] ^ d[237] ^ d[236] ^ d[235] ^ d[233] ^ d[232] ^ d[228] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[221] ^ d[217] ^ d[216] ^ d[214] ^ d[212] ^ d[210] ^ d[207] ^ d[205] ^ d[204] ^ d[201] ^ d[198] ^ d[195] ^ d[194] ^ d[191] ^ d[190] ^ d[189] ^ d[188] ^ d[187] ^ d[186] ^ d[184] ^ d[179] ^ d[178] ^ d[175] ^ d[172] ^ d[165] ^ d[162] ^ d[161] ^ d[160] ^ d[158] ^ d[156] ^ d[150] ^ d[149] ^ d[148] ^ d[146] ^ d[145] ^ d[143] ^ d[141] ^ d[140] ^ d[139] ^ d[136] ^ d[133] ^ d[132] ^ d[129] ^ d[126] ^ d[125] ^ d[124] ^ d[123] ^ d[121] ^ d[120] ^ d[117] ^ d[116] ^ d[115] ^ d[114] ^ d[110] ^ d[109] ^ d[108] ^ d[107] ^ d[105] ^ d[104] ^ d[102] ^ d[99] ^ d[96] ^ d[95] ^ d[94] ^ d[92] ^ d[91] ^ d[89] ^ d[88] ^ d[87] ^ d[83] ^ d[82] ^ d[80] ^ d[73] ^ d[71] ^ d[62] ^ d[61] ^ d[56] ^ d[53] ^ d[52] ^ d[51] ^ d[49] ^ d[42] ^ d[40] ^ d[37] ^ d[35] ^ d[34] ^ d[31] ^ d[29] ^ d[27] ^ d[26] ^ d[24] ^ d[22] ^ d[18] ^ d[17] ^ d[13] ^ d[10] ^ d[9] ^ d[5] ^ c[0] ^ c[4] ^ c[7] ^ c[8] ^ c[11] ^ c[14] ^ c[18] ^ c[19] ^ c[20] ^ c[21] ^ c[22] ^ c[24] ^ c[26] ^ c[27] ^ c[29] ^ c[30] ^ c[31];
    stage_2_crc_value[22] = d[506] ^ d[505] ^ d[503] ^ d[499] ^ d[494] ^ d[493] ^ d[491] ^ d[490] ^ d[486] ^ d[485] ^ d[483] ^ d[482] ^ d[479] ^ d[478] ^ d[477] ^ d[476] ^ d[470] ^ d[468] ^ d[463] ^ d[462] ^ d[460] ^ d[455] ^ d[452] ^ d[449] ^ d[448] ^ d[447] ^ d[446] ^ d[445] ^ d[444] ^ d[443] ^ d[442] ^ d[439] ^ d[438] ^ d[436] ^ d[435] ^ d[434] ^ d[430] ^ d[429] ^ d[427] ^ d[426] ^ d[424] ^ d[421] ^ d[420] ^ d[417] ^ d[413] ^ d[411] ^ d[410] ^ d[409] ^ d[408] ^ d[407] ^ d[405] ^ d[404] ^ d[402] ^ d[401] ^ d[400] ^ d[396] ^ d[395] ^ d[391] ^ d[389] ^ d[386] ^ d[385] ^ d[384] ^ d[381] ^ d[378] ^ d[377] ^ d[376] ^ d[375] ^ d[374] ^ d[373] ^ d[372] ^ d[370] ^ d[368] ^ d[367] ^ d[366] ^ d[362] ^ d[361] ^ d[358] ^ d[357] ^ d[355] ^ d[354] ^ d[346] ^ d[345] ^ d[343] ^ d[339] ^ d[338] ^ d[337] ^ d[336] ^ d[334] ^ d[330] ^ d[328] ^ d[326] ^ d[325] ^ d[321] ^ d[320] ^ d[319] ^ d[318] ^ d[317] ^ d[315] ^ d[313] ^ d[312] ^ d[311] ^ d[310] ^ d[308] ^ d[307] ^ d[306] ^ d[304] ^ d[300] ^ d[299] ^ d[297] ^ d[295] ^ d[293] ^ d[286] ^ d[283] ^ d[282] ^ d[280] ^ d[279] ^ d[277] ^ d[273] ^ d[270] ^ d[268] ^ d[266] ^ d[265] ^ d[264] ^ d[261] ^ d[259] ^ d[257] ^ d[256] ^ d[253] ^ d[251] ^ d[249] ^ d[248] ^ d[245] ^ d[244] ^ d[239] ^ d[238] ^ d[236] ^ d[233] ^ d[230] ^ d[229] ^ d[225] ^ d[222] ^ d[218] ^ d[217] ^ d[216] ^ d[215] ^ d[214] ^ d[213] ^ d[212] ^ d[211] ^ d[210] ^ d[209] ^ d[207] ^ d[206] ^ d[205] ^ d[203] ^ d[201] ^ d[198] ^ d[197] ^ d[196] ^ d[195] ^ d[194] ^ d[193] ^ d[189] ^ d[187] ^ d[186] ^ d[185] ^ d[183] ^ d[182] ^ d[180] ^ d[179] ^ d[176] ^ d[173] ^ d[172] ^ d[171] ^ d[170] ^ d[169] ^ d[167] ^ d[163] ^ d[159] ^ d[158] ^ d[157] ^ d[156] ^ d[155] ^ d[150] ^ d[147] ^ d[146] ^ d[143] ^ d[142] ^ d[141] ^ d[140] ^ d[136] ^ d[135] ^ d[133] ^ d[132] ^ d[130] ^ d[128] ^ d[124] ^ d[123] ^ d[122] ^ d[121] ^ d[119] ^ d[115] ^ d[114] ^ d[113] ^ d[109] ^ d[108] ^ d[105] ^ d[104] ^ d[101] ^ d[100] ^ d[99] ^ d[98] ^ d[94] ^ d[93] ^ d[92] ^ d[90] ^ d[89] ^ d[88] ^ d[87] ^ d[85] ^ d[82] ^ d[79] ^ d[74] ^ d[73] ^ d[68] ^ d[67] ^ d[66] ^ d[65] ^ d[62] ^ d[61] ^ d[60] ^ d[58] ^ d[57] ^ d[55] ^ d[52] ^ d[48] ^ d[47] ^ d[45] ^ d[44] ^ d[43] ^ d[41] ^ d[38] ^ d[37] ^ d[36] ^ d[35] ^ d[34] ^ d[31] ^ d[29] ^ d[27] ^ d[26] ^ d[24] ^ d[23] ^ d[19] ^ d[18] ^ d[16] ^ d[14] ^ d[12] ^ d[11] ^ d[9] ^ d[0] ^ c[2] ^ c[3] ^ c[5] ^ c[6] ^ c[10] ^ c[11] ^ c[13] ^ c[14] ^ c[19] ^ c[23] ^ c[25] ^ c[26];
    stage_2_crc_value[23] = d[511] ^ d[510] ^ d[508] ^ d[504] ^ d[502] ^ d[501] ^ d[493] ^ d[490] ^ d[489] ^ d[488] ^ d[487] ^ d[484] ^ d[482] ^ d[481] ^ d[478] ^ d[476] ^ d[472] ^ d[471] ^ d[470] ^ d[469] ^ d[468] ^ d[465] ^ d[463] ^ d[462] ^ d[458] ^ d[456] ^ d[453] ^ d[452] ^ d[447] ^ d[446] ^ d[445] ^ d[443] ^ d[440] ^ d[439] ^ d[435] ^ d[434] ^ d[433] ^ d[431] ^ d[430] ^ d[428] ^ d[427] ^ d[425] ^ d[424] ^ d[421] ^ d[419] ^ d[416] ^ d[411] ^ d[410] ^ d[407] ^ d[406] ^ d[404] ^ d[403] ^ d[402] ^ d[401] ^ d[400] ^ d[399] ^ d[398] ^ d[397] ^ d[393] ^ d[391] ^ d[388] ^ d[385] ^ d[382] ^ d[381] ^ d[379] ^ d[377] ^ d[375] ^ d[373] ^ d[372] ^ d[371] ^ d[367] ^ d[366] ^ d[357] ^ d[356] ^ d[355] ^ d[353] ^ d[349] ^ d[348] ^ d[346] ^ d[345] ^ d[342] ^ d[341] ^ d[340] ^ d[334] ^ d[333] ^ d[331] ^ d[329] ^ d[328] ^ d[326] ^ d[317] ^ d[316] ^ d[315] ^ d[314] ^ d[313] ^ d[311] ^ d[310] ^ d[308] ^ d[307] ^ d[303] ^ d[302] ^ d[301] ^ d[299] ^ d[297] ^ d[295] ^ d[292] ^ d[290] ^ d[288] ^ d[286] ^ d[284] ^ d[281] ^ d[280] ^ d[279] ^ d[278] ^ d[277] ^ d[276] ^ d[273] ^ d[271] ^ d[268] ^ d[267] ^ d[266] ^ d[264] ^ d[262] ^ d[261] ^ d[260] ^ d[259] ^ d[258] ^ d[255] ^ d[254] ^ d[250] ^ d[249] ^ d[248] ^ d[246] ^ d[245] ^ d[243] ^ d[240] ^ d[239] ^ d[231] ^ d[228] ^ d[227] ^ d[224] ^ d[223] ^ d[219] ^ d[218] ^ d[217] ^ d[215] ^ d[213] ^ d[211] ^ d[209] ^ d[206] ^ d[204] ^ d[203] ^ d[201] ^ d[196] ^ d[195] ^ d[193] ^ d[192] ^ d[191] ^ d[187] ^ d[184] ^ d[182] ^ d[181] ^ d[180] ^ d[177] ^ d[174] ^ d[173] ^ d[169] ^ d[168] ^ d[167] ^ d[166] ^ d[164] ^ d[162] ^ d[161] ^ d[160] ^ d[159] ^ d[157] ^ d[155] ^ d[149] ^ d[148] ^ d[147] ^ d[142] ^ d[141] ^ d[135] ^ d[133] ^ d[132] ^ d[131] ^ d[129] ^ d[128] ^ d[127] ^ d[126] ^ d[124] ^ d[122] ^ d[120] ^ d[119] ^ d[118] ^ d[117] ^ d[115] ^ d[113] ^ d[111] ^ d[109] ^ d[105] ^ d[104] ^ d[103] ^ d[102] ^ d[100] ^ d[98] ^ d[97] ^ d[96] ^ d[93] ^ d[91] ^ d[90] ^ d[89] ^ d[88] ^ d[87] ^ d[86] ^ d[85] ^ d[84] ^ d[82] ^ d[81] ^ d[80] ^ d[79] ^ d[75] ^ d[74] ^ d[73] ^ d[72] ^ d[69] ^ d[65] ^ d[62] ^ d[60] ^ d[59] ^ d[56] ^ d[55] ^ d[54] ^ d[50] ^ d[49] ^ d[47] ^ d[46] ^ d[42] ^ d[39] ^ d[38] ^ d[36] ^ d[35] ^ d[34] ^ d[31] ^ d[29] ^ d[27] ^ d[26] ^ d[20] ^ d[19] ^ d[17] ^ d[16] ^ d[15] ^ d[13] ^ d[9] ^ d[6] ^ d[1] ^ d[0] ^ c[1] ^ c[2] ^ c[4] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[13] ^ c[21] ^ c[22] ^ c[24] ^ c[28] ^ c[30] ^ c[31];
    stage_2_crc_value[24] = d[511] ^ d[509] ^ d[505] ^ d[503] ^ d[502] ^ d[494] ^ d[491] ^ d[490] ^ d[489] ^ d[488] ^ d[485] ^ d[483] ^ d[482] ^ d[479] ^ d[477] ^ d[473] ^ d[472] ^ d[471] ^ d[470] ^ d[469] ^ d[466] ^ d[464] ^ d[463] ^ d[459] ^ d[457] ^ d[454] ^ d[453] ^ d[448] ^ d[447] ^ d[446] ^ d[444] ^ d[441] ^ d[440] ^ d[436] ^ d[435] ^ d[434] ^ d[432] ^ d[431] ^ d[429] ^ d[428] ^ d[426] ^ d[425] ^ d[422] ^ d[420] ^ d[417] ^ d[412] ^ d[411] ^ d[408] ^ d[407] ^ d[405] ^ d[404] ^ d[403] ^ d[402] ^ d[401] ^ d[400] ^ d[399] ^ d[398] ^ d[394] ^ d[392] ^ d[389] ^ d[386] ^ d[383] ^ d[382] ^ d[380] ^ d[378] ^ d[376] ^ d[374] ^ d[373] ^ d[372] ^ d[368] ^ d[367] ^ d[358] ^ d[357] ^ d[356] ^ d[354] ^ d[350] ^ d[349] ^ d[347] ^ d[346] ^ d[343] ^ d[342] ^ d[341] ^ d[335] ^ d[334] ^ d[332] ^ d[330] ^ d[329] ^ d[327] ^ d[318] ^ d[317] ^ d[316] ^ d[315] ^ d[314] ^ d[312] ^ d[311] ^ d[309] ^ d[308] ^ d[304] ^ d[303] ^ d[302] ^ d[300] ^ d[298] ^ d[296] ^ d[293] ^ d[291] ^ d[289] ^ d[287] ^ d[285] ^ d[282] ^ d[281] ^ d[280] ^ d[279] ^ d[278] ^ d[277] ^ d[274] ^ d[272] ^ d[269] ^ d[268] ^ d[267] ^ d[265] ^ d[263] ^ d[262] ^ d[261] ^ d[260] ^ d[259] ^ d[256] ^ d[255] ^ d[251] ^ d[250] ^ d[249] ^ d[247] ^ d[246] ^ d[244] ^ d[241] ^ d[240] ^ d[232] ^ d[229] ^ d[228] ^ d[225] ^ d[224] ^ d[220] ^ d[219] ^ d[218] ^ d[216] ^ d[214] ^ d[212] ^ d[210] ^ d[207] ^ d[205] ^ d[204] ^ d[202] ^ d[197] ^ d[196] ^ d[194] ^ d[193] ^ d[192] ^ d[188] ^ d[185] ^ d[183] ^ d[182] ^ d[181] ^ d[178] ^ d[175] ^ d[174] ^ d[170] ^ d[169] ^ d[168] ^ d[167] ^ d[165] ^ d[163] ^ d[162] ^ d[161] ^ d[160] ^ d[158] ^ d[156] ^ d[150] ^ d[149] ^ d[148] ^ d[143] ^ d[142] ^ d[136] ^ d[134] ^ d[133] ^ d[132] ^ d[130] ^ d[129] ^ d[128] ^ d[127] ^ d[125] ^ d[123] ^ d[121] ^ d[120] ^ d[119] ^ d[118] ^ d[116] ^ d[114] ^ d[112] ^ d[110] ^ d[106] ^ d[105] ^ d[104] ^ d[103] ^ d[101] ^ d[99] ^ d[98] ^ d[97] ^ d[94] ^ d[92] ^ d[91] ^ d[90] ^ d[89] ^ d[88] ^ d[87] ^ d[86] ^ d[85] ^ d[83] ^ d[82] ^ d[81] ^ d[80] ^ d[76] ^ d[75] ^ d[74] ^ d[73] ^ d[70] ^ d[66] ^ d[63] ^ d[61] ^ d[60] ^ d[57] ^ d[56] ^ d[55] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[43] ^ d[40] ^ d[39] ^ d[37] ^ d[36] ^ d[35] ^ d[32] ^ d[30] ^ d[28] ^ d[27] ^ d[21] ^ d[20] ^ d[18] ^ d[17] ^ d[16] ^ d[14] ^ d[10] ^ d[7] ^ d[2] ^ d[1] ^ c[2] ^ c[3] ^ c[5] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[14] ^ c[22] ^ c[23] ^ c[25] ^ c[29] ^ c[31];
    stage_2_crc_value[25] = d[510] ^ d[506] ^ d[504] ^ d[503] ^ d[495] ^ d[492] ^ d[491] ^ d[490] ^ d[489] ^ d[486] ^ d[484] ^ d[483] ^ d[480] ^ d[478] ^ d[474] ^ d[473] ^ d[472] ^ d[471] ^ d[470] ^ d[467] ^ d[465] ^ d[464] ^ d[460] ^ d[458] ^ d[455] ^ d[454] ^ d[449] ^ d[448] ^ d[447] ^ d[445] ^ d[442] ^ d[441] ^ d[437] ^ d[436] ^ d[435] ^ d[433] ^ d[432] ^ d[430] ^ d[429] ^ d[427] ^ d[426] ^ d[423] ^ d[421] ^ d[418] ^ d[413] ^ d[412] ^ d[409] ^ d[408] ^ d[406] ^ d[405] ^ d[404] ^ d[403] ^ d[402] ^ d[401] ^ d[400] ^ d[399] ^ d[395] ^ d[393] ^ d[390] ^ d[387] ^ d[384] ^ d[383] ^ d[381] ^ d[379] ^ d[377] ^ d[375] ^ d[374] ^ d[373] ^ d[369] ^ d[368] ^ d[359] ^ d[358] ^ d[357] ^ d[355] ^ d[351] ^ d[350] ^ d[348] ^ d[347] ^ d[344] ^ d[343] ^ d[342] ^ d[336] ^ d[335] ^ d[333] ^ d[331] ^ d[330] ^ d[328] ^ d[319] ^ d[318] ^ d[317] ^ d[316] ^ d[315] ^ d[313] ^ d[312] ^ d[310] ^ d[309] ^ d[305] ^ d[304] ^ d[303] ^ d[301] ^ d[299] ^ d[297] ^ d[294] ^ d[292] ^ d[290] ^ d[288] ^ d[286] ^ d[283] ^ d[282] ^ d[281] ^ d[280] ^ d[279] ^ d[278] ^ d[275] ^ d[273] ^ d[270] ^ d[269] ^ d[268] ^ d[266] ^ d[264] ^ d[263] ^ d[262] ^ d[261] ^ d[260] ^ d[257] ^ d[256] ^ d[252] ^ d[251] ^ d[250] ^ d[248] ^ d[247] ^ d[245] ^ d[242] ^ d[241] ^ d[233] ^ d[230] ^ d[229] ^ d[226] ^ d[225] ^ d[221] ^ d[220] ^ d[219] ^ d[217] ^ d[215] ^ d[213] ^ d[211] ^ d[208] ^ d[206] ^ d[205] ^ d[203] ^ d[198] ^ d[197] ^ d[195] ^ d[194] ^ d[193] ^ d[189] ^ d[186] ^ d[184] ^ d[183] ^ d[182] ^ d[179] ^ d[176] ^ d[175] ^ d[171] ^ d[170] ^ d[169] ^ d[168] ^ d[166] ^ d[164] ^ d[163] ^ d[162] ^ d[161] ^ d[159] ^ d[157] ^ d[151] ^ d[150] ^ d[149] ^ d[144] ^ d[143] ^ d[137] ^ d[135] ^ d[134] ^ d[133] ^ d[131] ^ d[130] ^ d[129] ^ d[128] ^ d[126] ^ d[124] ^ d[122] ^ d[121] ^ d[120] ^ d[119] ^ d[117] ^ d[115] ^ d[113] ^ d[111] ^ d[107] ^ d[106] ^ d[105] ^ d[104] ^ d[102] ^ d[100] ^ d[99] ^ d[98] ^ d[95] ^ d[93] ^ d[92] ^ d[91] ^ d[90] ^ d[89] ^ d[88] ^ d[87] ^ d[86] ^ d[84] ^ d[83] ^ d[82] ^ d[81] ^ d[77] ^ d[76] ^ d[75] ^ d[74] ^ d[71] ^ d[67] ^ d[64] ^ d[62] ^ d[61] ^ d[58] ^ d[57] ^ d[56] ^ d[52] ^ d[51] ^ d[49] ^ d[48] ^ d[44] ^ d[41] ^ d[40] ^ d[38] ^ d[37] ^ d[36] ^ d[33] ^ d[31] ^ d[29] ^ d[28] ^ d[22] ^ d[21] ^ d[19] ^ d[18] ^ d[17] ^ d[15] ^ d[11] ^ d[8] ^ d[3] ^ d[2] ^ c[0] ^ c[3] ^ c[4] ^ c[6] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[15] ^ c[23] ^ c[24] ^ c[26] ^ c[30];
    stage_2_crc_value[26] = d[510] ^ d[508] ^ d[506] ^ d[505] ^ d[504] ^ d[502] ^ d[501] ^ d[500] ^ d[496] ^ d[495] ^ d[494] ^ d[489] ^ d[488] ^ d[487] ^ d[486] ^ d[485] ^ d[484] ^ d[483] ^ d[482] ^ d[480] ^ d[477] ^ d[476] ^ d[475] ^ d[474] ^ d[473] ^ d[471] ^ d[470] ^ d[466] ^ d[464] ^ d[462] ^ d[459] ^ d[458] ^ d[456] ^ d[455] ^ d[452] ^ d[446] ^ d[444] ^ d[443] ^ d[442] ^ d[438] ^ d[431] ^ d[430] ^ d[428] ^ d[427] ^ d[418] ^ d[416] ^ d[413] ^ d[412] ^ d[410] ^ d[408] ^ d[406] ^ d[403] ^ d[402] ^ d[401] ^ d[399] ^ d[398] ^ d[394] ^ d[393] ^ d[392] ^ d[390] ^ d[387] ^ d[386] ^ d[385] ^ d[384] ^ d[382] ^ d[381] ^ d[380] ^ d[375] ^ d[372] ^ d[370] ^ d[368] ^ d[366] ^ d[363] ^ d[362] ^ d[360] ^ d[357] ^ d[356] ^ d[353] ^ d[352] ^ d[351] ^ d[347] ^ d[343] ^ d[342] ^ d[341] ^ d[339] ^ d[338] ^ d[336] ^ d[335] ^ d[333] ^ d[332] ^ d[331] ^ d[329] ^ d[328] ^ d[327] ^ d[322] ^ d[321] ^ d[316] ^ d[315] ^ d[314] ^ d[313] ^ d[312] ^ d[311] ^ d[309] ^ d[306] ^ d[304] ^ d[303] ^ d[299] ^ d[297] ^ d[296] ^ d[294] ^ d[293] ^ d[292] ^ d[291] ^ d[290] ^ d[289] ^ d[288] ^ d[286] ^ d[284] ^ d[282] ^ d[281] ^ d[280] ^ d[277] ^ d[273] ^ d[271] ^ d[270] ^ d[268] ^ d[267] ^ d[263] ^ d[262] ^ d[259] ^ d[258] ^ d[255] ^ d[253] ^ d[251] ^ d[249] ^ d[246] ^ d[242] ^ d[237] ^ d[231] ^ d[228] ^ d[224] ^ d[222] ^ d[221] ^ d[220] ^ d[218] ^ d[210] ^ d[208] ^ d[206] ^ d[204] ^ d[203] ^ d[202] ^ d[201] ^ d[197] ^ d[196] ^ d[195] ^ d[193] ^ d[192] ^ d[191] ^ d[188] ^ d[187] ^ d[186] ^ d[185] ^ d[184] ^ d[182] ^ d[180] ^ d[177] ^ d[176] ^ d[166] ^ d[165] ^ d[164] ^ d[163] ^ d[161] ^ d[160] ^ d[156] ^ d[155] ^ d[152] ^ d[150] ^ d[149] ^ d[145] ^ d[143] ^ d[138] ^ d[137] ^ d[131] ^ d[130] ^ d[129] ^ d[128] ^ d[126] ^ d[122] ^ d[121] ^ d[120] ^ d[119] ^ d[117] ^ d[113] ^ d[112] ^ d[111] ^ d[110] ^ d[108] ^ d[107] ^ d[105] ^ d[104] ^ d[100] ^ d[98] ^ d[97] ^ d[95] ^ d[93] ^ d[92] ^ d[91] ^ d[90] ^ d[89] ^ d[88] ^ d[81] ^ d[79] ^ d[78] ^ d[77] ^ d[76] ^ d[75] ^ d[73] ^ d[67] ^ d[66] ^ d[62] ^ d[61] ^ d[60] ^ d[59] ^ d[57] ^ d[55] ^ d[54] ^ d[52] ^ d[49] ^ d[48] ^ d[47] ^ d[44] ^ d[42] ^ d[41] ^ d[39] ^ d[38] ^ d[31] ^ d[28] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[20] ^ d[19] ^ d[18] ^ d[10] ^ d[6] ^ d[4] ^ d[3] ^ d[0] ^ c[0] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[14] ^ c[15] ^ c[16] ^ c[20] ^ c[21] ^ c[22] ^ c[24] ^ c[25] ^ c[26] ^ c[28] ^ c[30];
    stage_2_crc_value[27] = d[511] ^ d[509] ^ d[507] ^ d[506] ^ d[505] ^ d[503] ^ d[502] ^ d[501] ^ d[497] ^ d[496] ^ d[495] ^ d[490] ^ d[489] ^ d[488] ^ d[487] ^ d[486] ^ d[485] ^ d[484] ^ d[483] ^ d[481] ^ d[478] ^ d[477] ^ d[476] ^ d[475] ^ d[474] ^ d[472] ^ d[471] ^ d[467] ^ d[465] ^ d[463] ^ d[460] ^ d[459] ^ d[457] ^ d[456] ^ d[453] ^ d[447] ^ d[445] ^ d[444] ^ d[443] ^ d[439] ^ d[432] ^ d[431] ^ d[429] ^ d[428] ^ d[419] ^ d[417] ^ d[414] ^ d[413] ^ d[411] ^ d[409] ^ d[407] ^ d[404] ^ d[403] ^ d[402] ^ d[400] ^ d[399] ^ d[395] ^ d[394] ^ d[393] ^ d[391] ^ d[388] ^ d[387] ^ d[386] ^ d[385] ^ d[383] ^ d[382] ^ d[381] ^ d[376] ^ d[373] ^ d[371] ^ d[369] ^ d[367] ^ d[364] ^ d[363] ^ d[361] ^ d[358] ^ d[357] ^ d[354] ^ d[353] ^ d[352] ^ d[348] ^ d[344] ^ d[343] ^ d[342] ^ d[340] ^ d[339] ^ d[337] ^ d[336] ^ d[334] ^ d[333] ^ d[332] ^ d[330] ^ d[329] ^ d[328] ^ d[323] ^ d[322] ^ d[317] ^ d[316] ^ d[315] ^ d[314] ^ d[313] ^ d[312] ^ d[310] ^ d[307] ^ d[305] ^ d[304] ^ d[300] ^ d[298] ^ d[297] ^ d[295] ^ d[294] ^ d[293] ^ d[292] ^ d[291] ^ d[290] ^ d[289] ^ d[287] ^ d[285] ^ d[283] ^ d[282] ^ d[281] ^ d[278] ^ d[274] ^ d[272] ^ d[271] ^ d[269] ^ d[268] ^ d[264] ^ d[263] ^ d[260] ^ d[259] ^ d[256] ^ d[254] ^ d[252] ^ d[250] ^ d[247] ^ d[243] ^ d[238] ^ d[232] ^ d[229] ^ d[225] ^ d[223] ^ d[222] ^ d[221] ^ d[219] ^ d[211] ^ d[209] ^ d[207] ^ d[205] ^ d[204] ^ d[203] ^ d[202] ^ d[198] ^ d[197] ^ d[196] ^ d[194] ^ d[193] ^ d[192] ^ d[189] ^ d[188] ^ d[187] ^ d[186] ^ d[185] ^ d[183] ^ d[181] ^ d[178] ^ d[177] ^ d[167] ^ d[166] ^ d[165] ^ d[164] ^ d[162] ^ d[161] ^ d[157] ^ d[156] ^ d[153] ^ d[151] ^ d[150] ^ d[146] ^ d[144] ^ d[139] ^ d[138] ^ d[132] ^ d[131] ^ d[130] ^ d[129] ^ d[127] ^ d[123] ^ d[122] ^ d[121] ^ d[120] ^ d[118] ^ d[114] ^ d[113] ^ d[112] ^ d[111] ^ d[109] ^ d[108] ^ d[106] ^ d[105] ^ d[101] ^ d[99] ^ d[98] ^ d[96] ^ d[94] ^ d[93] ^ d[92] ^ d[91] ^ d[90] ^ d[89] ^ d[82] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[76] ^ d[74] ^ d[68] ^ d[67] ^ d[63] ^ d[62] ^ d[61] ^ d[60] ^ d[58] ^ d[56] ^ d[55] ^ d[53] ^ d[50] ^ d[49] ^ d[48] ^ d[45] ^ d[43] ^ d[42] ^ d[40] ^ d[39] ^ d[32] ^ d[29] ^ d[27] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[21] ^ d[20] ^ d[19] ^ d[11] ^ d[7] ^ d[5] ^ d[4] ^ d[1] ^ c[1] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[15] ^ c[16] ^ c[17] ^ c[21] ^ c[22] ^ c[23] ^ c[25] ^ c[26] ^ c[27] ^ c[29] ^ c[31];
    stage_2_crc_value[28] = d[510] ^ d[508] ^ d[507] ^ d[506] ^ d[504] ^ d[503] ^ d[502] ^ d[498] ^ d[497] ^ d[496] ^ d[491] ^ d[490] ^ d[489] ^ d[488] ^ d[487] ^ d[486] ^ d[485] ^ d[484] ^ d[482] ^ d[479] ^ d[478] ^ d[477] ^ d[476] ^ d[475] ^ d[473] ^ d[472] ^ d[468] ^ d[466] ^ d[464] ^ d[461] ^ d[460] ^ d[458] ^ d[457] ^ d[454] ^ d[448] ^ d[446] ^ d[445] ^ d[444] ^ d[440] ^ d[433] ^ d[432] ^ d[430] ^ d[429] ^ d[420] ^ d[418] ^ d[415] ^ d[414] ^ d[412] ^ d[410] ^ d[408] ^ d[405] ^ d[404] ^ d[403] ^ d[401] ^ d[400] ^ d[396] ^ d[395] ^ d[394] ^ d[392] ^ d[389] ^ d[388] ^ d[387] ^ d[386] ^ d[384] ^ d[383] ^ d[382] ^ d[377] ^ d[374] ^ d[372] ^ d[370] ^ d[368] ^ d[365] ^ d[364] ^ d[362] ^ d[359] ^ d[358] ^ d[355] ^ d[354] ^ d[353] ^ d[349] ^ d[345] ^ d[344] ^ d[343] ^ d[341] ^ d[340] ^ d[338] ^ d[337] ^ d[335] ^ d[334] ^ d[333] ^ d[331] ^ d[330] ^ d[329] ^ d[324] ^ d[323] ^ d[318] ^ d[317] ^ d[316] ^ d[315] ^ d[314] ^ d[313] ^ d[311] ^ d[308] ^ d[306] ^ d[305] ^ d[301] ^ d[299] ^ d[298] ^ d[296] ^ d[295] ^ d[294] ^ d[293] ^ d[292] ^ d[291] ^ d[290] ^ d[288] ^ d[286] ^ d[284] ^ d[283] ^ d[282] ^ d[279] ^ d[275] ^ d[273] ^ d[272] ^ d[270] ^ d[269] ^ d[265] ^ d[264] ^ d[261] ^ d[260] ^ d[257] ^ d[255] ^ d[253] ^ d[251] ^ d[248] ^ d[244] ^ d[239] ^ d[233] ^ d[230] ^ d[226] ^ d[224] ^ d[223] ^ d[222] ^ d[220] ^ d[212] ^ d[210] ^ d[208] ^ d[206] ^ d[205] ^ d[204] ^ d[203] ^ d[199] ^ d[198] ^ d[197] ^ d[195] ^ d[194] ^ d[193] ^ d[190] ^ d[189] ^ d[188] ^ d[187] ^ d[186] ^ d[184] ^ d[182] ^ d[179] ^ d[178] ^ d[168] ^ d[167] ^ d[166] ^ d[165] ^ d[163] ^ d[162] ^ d[158] ^ d[157] ^ d[154] ^ d[152] ^ d[151] ^ d[147] ^ d[145] ^ d[140] ^ d[139] ^ d[133] ^ d[132] ^ d[131] ^ d[130] ^ d[128] ^ d[124] ^ d[123] ^ d[122] ^ d[121] ^ d[119] ^ d[115] ^ d[114] ^ d[113] ^ d[112] ^ d[110] ^ d[109] ^ d[107] ^ d[106] ^ d[102] ^ d[100] ^ d[99] ^ d[97] ^ d[95] ^ d[94] ^ d[93] ^ d[92] ^ d[91] ^ d[90] ^ d[83] ^ d[81] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[75] ^ d[69] ^ d[68] ^ d[64] ^ d[63] ^ d[62] ^ d[61] ^ d[59] ^ d[57] ^ d[56] ^ d[54] ^ d[51] ^ d[50] ^ d[49] ^ d[46] ^ d[44] ^ d[43] ^ d[41] ^ d[40] ^ d[33] ^ d[30] ^ d[28] ^ d[27] ^ d[26] ^ d[25] ^ d[24] ^ d[22] ^ d[21] ^ d[20] ^ d[12] ^ d[8] ^ d[6] ^ d[5] ^ d[2] ^ c[2] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[16] ^ c[17] ^ c[18] ^ c[22] ^ c[23] ^ c[24] ^ c[26] ^ c[27] ^ c[28] ^ c[30];
    stage_2_crc_value[29] = d[511] ^ d[509] ^ d[508] ^ d[507] ^ d[505] ^ d[504] ^ d[503] ^ d[499] ^ d[498] ^ d[497] ^ d[492] ^ d[491] ^ d[490] ^ d[489] ^ d[488] ^ d[487] ^ d[486] ^ d[485] ^ d[483] ^ d[480] ^ d[479] ^ d[478] ^ d[477] ^ d[476] ^ d[474] ^ d[473] ^ d[469] ^ d[467] ^ d[465] ^ d[462] ^ d[461] ^ d[459] ^ d[458] ^ d[455] ^ d[449] ^ d[447] ^ d[446] ^ d[445] ^ d[441] ^ d[434] ^ d[433] ^ d[431] ^ d[430] ^ d[421] ^ d[419] ^ d[416] ^ d[415] ^ d[413] ^ d[411] ^ d[409] ^ d[406] ^ d[405] ^ d[404] ^ d[402] ^ d[401] ^ d[397] ^ d[396] ^ d[395] ^ d[393] ^ d[390] ^ d[389] ^ d[388] ^ d[387] ^ d[385] ^ d[384] ^ d[383] ^ d[378] ^ d[375] ^ d[373] ^ d[371] ^ d[369] ^ d[366] ^ d[365] ^ d[363] ^ d[360] ^ d[359] ^ d[356] ^ d[355] ^ d[354] ^ d[350] ^ d[346] ^ d[345] ^ d[344] ^ d[342] ^ d[341] ^ d[339] ^ d[338] ^ d[336] ^ d[335] ^ d[334] ^ d[332] ^ d[331] ^ d[330] ^ d[325] ^ d[324] ^ d[319] ^ d[318] ^ d[317] ^ d[316] ^ d[315] ^ d[314] ^ d[312] ^ d[309] ^ d[307] ^ d[306] ^ d[302] ^ d[300] ^ d[299] ^ d[297] ^ d[296] ^ d[295] ^ d[294] ^ d[293] ^ d[292] ^ d[291] ^ d[289] ^ d[287] ^ d[285] ^ d[284] ^ d[283] ^ d[280] ^ d[276] ^ d[274] ^ d[273] ^ d[271] ^ d[270] ^ d[266] ^ d[265] ^ d[262] ^ d[261] ^ d[258] ^ d[256] ^ d[254] ^ d[252] ^ d[249] ^ d[245] ^ d[240] ^ d[234] ^ d[231] ^ d[227] ^ d[225] ^ d[224] ^ d[223] ^ d[221] ^ d[213] ^ d[211] ^ d[209] ^ d[207] ^ d[206] ^ d[205] ^ d[204] ^ d[200] ^ d[199] ^ d[198] ^ d[196] ^ d[195] ^ d[194] ^ d[191] ^ d[190] ^ d[189] ^ d[188] ^ d[187] ^ d[185] ^ d[183] ^ d[180] ^ d[179] ^ d[169] ^ d[168] ^ d[167] ^ d[166] ^ d[164] ^ d[163] ^ d[159] ^ d[158] ^ d[155] ^ d[153] ^ d[152] ^ d[148] ^ d[146] ^ d[141] ^ d[140] ^ d[134] ^ d[133] ^ d[132] ^ d[131] ^ d[129] ^ d[125] ^ d[124] ^ d[123] ^ d[122] ^ d[120] ^ d[116] ^ d[115] ^ d[114] ^ d[113] ^ d[111] ^ d[110] ^ d[108] ^ d[107] ^ d[103] ^ d[101] ^ d[100] ^ d[98] ^ d[96] ^ d[95] ^ d[94] ^ d[93] ^ d[92] ^ d[91] ^ d[84] ^ d[82] ^ d[81] ^ d[80] ^ d[79] ^ d[78] ^ d[76] ^ d[70] ^ d[69] ^ d[65] ^ d[64] ^ d[63] ^ d[62] ^ d[60] ^ d[58] ^ d[57] ^ d[55] ^ d[52] ^ d[51] ^ d[50] ^ d[47] ^ d[45] ^ d[44] ^ d[42] ^ d[41] ^ d[34] ^ d[31] ^ d[29] ^ d[28] ^ d[27] ^ d[26] ^ d[25] ^ d[23] ^ d[22] ^ d[21] ^ d[13] ^ d[9] ^ d[7] ^ d[6] ^ d[3] ^ c[0] ^ c[3] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[17] ^ c[18] ^ c[19] ^ c[23] ^ c[24] ^ c[25] ^ c[27] ^ c[28] ^ c[29] ^ c[31];
    stage_2_crc_value[30] = d[510] ^ d[509] ^ d[508] ^ d[506] ^ d[505] ^ d[504] ^ d[500] ^ d[499] ^ d[498] ^ d[493] ^ d[492] ^ d[491] ^ d[490] ^ d[489] ^ d[488] ^ d[487] ^ d[486] ^ d[484] ^ d[481] ^ d[480] ^ d[479] ^ d[478] ^ d[477] ^ d[475] ^ d[474] ^ d[470] ^ d[468] ^ d[466] ^ d[463] ^ d[462] ^ d[460] ^ d[459] ^ d[456] ^ d[450] ^ d[448] ^ d[447] ^ d[446] ^ d[442] ^ d[435] ^ d[434] ^ d[432] ^ d[431] ^ d[422] ^ d[420] ^ d[417] ^ d[416] ^ d[414] ^ d[412] ^ d[410] ^ d[407] ^ d[406] ^ d[405] ^ d[403] ^ d[402] ^ d[398] ^ d[397] ^ d[396] ^ d[394] ^ d[391] ^ d[390] ^ d[389] ^ d[388] ^ d[386] ^ d[385] ^ d[384] ^ d[379] ^ d[376] ^ d[374] ^ d[372] ^ d[370] ^ d[367] ^ d[366] ^ d[364] ^ d[361] ^ d[360] ^ d[357] ^ d[356] ^ d[355] ^ d[351] ^ d[347] ^ d[346] ^ d[345] ^ d[343] ^ d[342] ^ d[340] ^ d[339] ^ d[337] ^ d[336] ^ d[335] ^ d[333] ^ d[332] ^ d[331] ^ d[326] ^ d[325] ^ d[320] ^ d[319] ^ d[318] ^ d[317] ^ d[316] ^ d[315] ^ d[313] ^ d[310] ^ d[308] ^ d[307] ^ d[303] ^ d[301] ^ d[300] ^ d[298] ^ d[297] ^ d[296] ^ d[295] ^ d[294] ^ d[293] ^ d[292] ^ d[290] ^ d[288] ^ d[286] ^ d[285] ^ d[284] ^ d[281] ^ d[277] ^ d[275] ^ d[274] ^ d[272] ^ d[271] ^ d[267] ^ d[266] ^ d[263] ^ d[262] ^ d[259] ^ d[257] ^ d[255] ^ d[253] ^ d[250] ^ d[246] ^ d[241] ^ d[235] ^ d[232] ^ d[228] ^ d[226] ^ d[225] ^ d[224] ^ d[222] ^ d[214] ^ d[212] ^ d[210] ^ d[208] ^ d[207] ^ d[206] ^ d[205] ^ d[201] ^ d[200] ^ d[199] ^ d[197] ^ d[196] ^ d[195] ^ d[192] ^ d[191] ^ d[190] ^ d[189] ^ d[188] ^ d[186] ^ d[184] ^ d[181] ^ d[180] ^ d[170] ^ d[169] ^ d[168] ^ d[167] ^ d[165] ^ d[164] ^ d[160] ^ d[159] ^ d[156] ^ d[154] ^ d[153] ^ d[149] ^ d[147] ^ d[142] ^ d[141] ^ d[135] ^ d[134] ^ d[133] ^ d[132] ^ d[130] ^ d[126] ^ d[125] ^ d[124] ^ d[123] ^ d[121] ^ d[117] ^ d[116] ^ d[115] ^ d[114] ^ d[112] ^ d[111] ^ d[109] ^ d[108] ^ d[104] ^ d[102] ^ d[101] ^ d[99] ^ d[97] ^ d[96] ^ d[95] ^ d[94] ^ d[93] ^ d[92] ^ d[85] ^ d[83] ^ d[82] ^ d[81] ^ d[80] ^ d[79] ^ d[77] ^ d[71] ^ d[70] ^ d[66] ^ d[65] ^ d[64] ^ d[63] ^ d[61] ^ d[59] ^ d[58] ^ d[56] ^ d[53] ^ d[52] ^ d[51] ^ d[48] ^ d[46] ^ d[45] ^ d[43] ^ d[42] ^ d[35] ^ d[32] ^ d[30] ^ d[29] ^ d[28] ^ d[27] ^ d[26] ^ d[24] ^ d[23] ^ d[22] ^ d[14] ^ d[10] ^ d[8] ^ d[7] ^ d[4] ^ c[0] ^ c[1] ^ c[4] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[18] ^ c[19] ^ c[20] ^ c[24] ^ c[25] ^ c[26] ^ c[28] ^ c[29] ^ c[30];
    stage_2_crc_value[31] = d[511] ^ d[510] ^ d[509] ^ d[507] ^ d[506] ^ d[505] ^ d[501] ^ d[500] ^ d[499] ^ d[494] ^ d[493] ^ d[492] ^ d[491] ^ d[490] ^ d[489] ^ d[488] ^ d[487] ^ d[485] ^ d[482] ^ d[481] ^ d[480] ^ d[479] ^ d[478] ^ d[476] ^ d[475] ^ d[471] ^ d[469] ^ d[467] ^ d[464] ^ d[463] ^ d[461] ^ d[460] ^ d[457] ^ d[451] ^ d[449] ^ d[448] ^ d[447] ^ d[443] ^ d[436] ^ d[435] ^ d[433] ^ d[432] ^ d[423] ^ d[421] ^ d[418] ^ d[417] ^ d[415] ^ d[413] ^ d[411] ^ d[408] ^ d[407] ^ d[406] ^ d[404] ^ d[403] ^ d[399] ^ d[398] ^ d[397] ^ d[395] ^ d[392] ^ d[391] ^ d[390] ^ d[389] ^ d[387] ^ d[386] ^ d[385] ^ d[380] ^ d[377] ^ d[375] ^ d[373] ^ d[371] ^ d[368] ^ d[367] ^ d[365] ^ d[362] ^ d[361] ^ d[358] ^ d[357] ^ d[356] ^ d[352] ^ d[348] ^ d[347] ^ d[346] ^ d[344] ^ d[343] ^ d[341] ^ d[340] ^ d[338] ^ d[337] ^ d[336] ^ d[334] ^ d[333] ^ d[332] ^ d[327] ^ d[326] ^ d[321] ^ d[320] ^ d[319] ^ d[318] ^ d[317] ^ d[316] ^ d[314] ^ d[311] ^ d[309] ^ d[308] ^ d[304] ^ d[302] ^ d[301] ^ d[299] ^ d[298] ^ d[297] ^ d[296] ^ d[295] ^ d[294] ^ d[293] ^ d[291] ^ d[289] ^ d[287] ^ d[286] ^ d[285] ^ d[282] ^ d[278] ^ d[276] ^ d[275] ^ d[273] ^ d[272] ^ d[268] ^ d[267] ^ d[264] ^ d[263] ^ d[260] ^ d[258] ^ d[256] ^ d[254] ^ d[251] ^ d[247] ^ d[242] ^ d[236] ^ d[233] ^ d[229] ^ d[227] ^ d[226] ^ d[225] ^ d[223] ^ d[215] ^ d[213] ^ d[211] ^ d[209] ^ d[208] ^ d[207] ^ d[206] ^ d[202] ^ d[201] ^ d[200] ^ d[198] ^ d[197] ^ d[196] ^ d[193] ^ d[192] ^ d[191] ^ d[190] ^ d[189] ^ d[187] ^ d[185] ^ d[182] ^ d[181] ^ d[171] ^ d[170] ^ d[169] ^ d[168] ^ d[166] ^ d[165] ^ d[161] ^ d[160] ^ d[157] ^ d[155] ^ d[154] ^ d[150] ^ d[148] ^ d[143] ^ d[142] ^ d[136] ^ d[135] ^ d[134] ^ d[133] ^ d[131] ^ d[127] ^ d[126] ^ d[125] ^ d[124] ^ d[122] ^ d[118] ^ d[117] ^ d[116] ^ d[115] ^ d[113] ^ d[112] ^ d[110] ^ d[109] ^ d[105] ^ d[103] ^ d[102] ^ d[100] ^ d[98] ^ d[97] ^ d[96] ^ d[95] ^ d[94] ^ d[93] ^ d[86] ^ d[84] ^ d[83] ^ d[82] ^ d[81] ^ d[80] ^ d[78] ^ d[72] ^ d[71] ^ d[67] ^ d[66] ^ d[65] ^ d[64] ^ d[62] ^ d[60] ^ d[59] ^ d[57] ^ d[54] ^ d[53] ^ d[52] ^ d[49] ^ d[47] ^ d[46] ^ d[44] ^ d[43] ^ d[36] ^ d[33] ^ d[31] ^ d[30] ^ d[29] ^ d[28] ^ d[27] ^ d[25] ^ d[24] ^ d[23] ^ d[15] ^ d[11] ^ d[9] ^ d[8] ^ d[5] ^ c[0] ^ c[1] ^ c[2] ^ c[5] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[19] ^ c[20] ^ c[21] ^ c[25] ^ c[26] ^ c[27] ^ c[29] ^ c[30] ^ c[31];

    
    ///////////////////////////////////////////////////////////////////////
    //
    // STAGE 3: CRC INSERTION
    //
    ///////////////////////////////////////////////////////////////////////
    
    // Forward direct values: 
    stage_3_valid <= stage_2_valid;
    stage_3_last <= stage_2_last;
    
    // Fill data word with bypassed value, CRC will be inserted later 
    stage_3_data <= stage_2_data_bypass; 

    // Insert the ICRC in the bypassed data - only applies if the current word is last
    if(stage_2_last) begin 
        // Based on keep, check if the word is full 
        if(stage_2_keep[63] == 1) begin
            stage_3_last <= 0; 
            stage_3_crc_value <= stage_2_crc_value; 
            // In this case, the pipeline must be stalled for one cycle to include the freshly formed word 
            stall_pipeline <= 1'b1; 
        end else begin 
            if(stage_2_last == 4'hf) begin
                stage_3_data[63:32] <= stage_2_crc_value; 
                stage_3_keep[7:4] <= 4'hf;
            end else if(stage_2_last == 8'hff) begin 
                stage_3_data[95:64] <= stage_2_crc_value; 
                stage_3_keep[11:8] <= 4'hf;
            end else if(stage_2_last == 12'hfff) begin 
                stage_3_data[127:96] <= stage_2_crc_value; 
                stage_3_keep[15:12] <= 4'hf;
            end else if(stage_2_last == 16'hffff) begin 
                stage_3_data[159:128] <= stage_2_crc_value; 
                stage_3_keep[19:16] <= 4'hf;
            end else if(stage_2_last == 20'hfffff) begin 
                stage_3_data[191:160] <= stage_2_crc_value; 
                stage_3_keep[23:20] <= 4'hf;
            end else if(stage_2_last == 24'hffffff) begin 
                stage_3_data[223:192] <= stage_2_crc_value; 
                stage_3_keep[27:24] <= 4'hf;
            end else if(stage_2_last == 28'hfffffff) begin
                stage_3_data[255:224] <= stage_2_crc_value; 
                stage_3_keep[31:28] <= 4'hf;
            end else if(stage_2_last == 32'hffffffff) begin 
                stage_3_data[287:256] <= stage_2_crc_value; 
                stage_3_keep[35:32] <= 4'hf;
            end else if(stage_2_last == 36'hfffffffff) begin
                stage_3_data[319:288] <= stage_2_crc_value; 
                stage_3_keep[39:36] <= 4'hf;
            end else if(stage_2_last == 40'hffffffffff) begin
                stage_3_data[351:320] <= stage_2_crc_value; 
                stage_3_keep[43:40] <= 4'hf;
            end else if(stage_2_last == 44'hfffffffffff) begin 
                stage_3_data[383:352] <= stage_2_crc_value; 
                stage_3_keep[47:44] <= 4'hf;
            end else if(stage_2_last == 48'hffffffffffff) begin 
                stage_3_data[415:384] <= stage_2_crc_value; 
                stage_3_keep[51:48] <= 4'hf;
            end else if(stage_2_last == 52'hfffffffffffff) begin
                stage_3_data[447:416] <= stage_2_crc_value; 
                stage_3_keep[55:52] <= 4'hf;
            end else if(stage_2_last == 56'hffffffffffffff) begin
                stage_3_data[479:448] <= stage_2_crc_value; 
                stage_3_keep[59:56] <= 4'hf;
            end else if(stage_2_last == 60'hfffffffffffffff) begin
                stage_3_data[511:480] <= stage_2_crc_value; 
                stage_3_keep[63:60] <= 4'hf;
            end
        end 

    end


    ///////////////////////////////////////////////////////////////////////
    //
    // STAGE 4: FORMATION OF A NEW WORD (if required)
    //
    ///////////////////////////////////////////////////////////////////////

    // Only act if pipeline is stalled 
    if(stall_pipeline) begin 
        switch_output <= 1; 
        stage_4_valid <= 1; 
        stage_4_last <= 1; 
        stage_4_data[31:0] <= stage_3_crc_value; 
        stage_4_data[511:32] <= 0; 
        stage_4_keep[3:0] <= 4'hf; 
        stage_4_keep[63:4] <= 0; 
        stall_pipeline <= 1'b0; 
    end else begin 
        switch_output <= 0; 
    end 
end 


//////////////////////////////////////////////////////////////////////////////////
//
// ASSIGN OUTPUTS TO THE PIPELINE
//
//////////////////////////////////////////////////////////////////////////////////

assign m_axis_tx.data = switch_output ? stage_4_data : stage_3_data; 
assign m_axis_tx.valid = switch_output ? stage_4_valid : stage_3_valid; 
assign m_axis_tx.last = switch_output ? stage_4_last : stage_3_last; 
assign m_axis_tx.keep = switch_output ? stage_4_keep : stage_3_keep; 


////////////////////////////////////////////////////////////////////////////////////
//
// ASSIGN READY INPUT TO THE PIPELINE
//
////////////////////////////////////////////////////////////////////////////////////

assign m_axis_rx.ready = m_axis_tx.ready; 




